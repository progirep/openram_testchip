VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project
  CLASS BLOCK ;
  FOREIGN user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 380.000 BY 414.000 ;
  PIN addrA0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 410.000 115.370 414.000 ;
    END
  END addrA0[0]
  PIN addrA0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END addrA0[1]
  PIN addrA0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END addrA0[2]
  PIN addrA0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END addrA0[3]
  PIN addrA0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END addrA0[4]
  PIN addrA0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END addrA0[5]
  PIN addrA0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END addrA0[6]
  PIN addrA0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END addrA0[7]
  PIN addrA1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 410.000 112.150 414.000 ;
    END
  END addrA1[0]
  PIN addrA1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 410.000 374.350 414.000 ;
    END
  END addrA1[1]
  PIN addrA1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 410.000 371.130 414.000 ;
    END
  END addrA1[2]
  PIN addrA1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 410.000 367.450 414.000 ;
    END
  END addrA1[3]
  PIN addrA1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 410.000 364.230 414.000 ;
    END
  END addrA1[4]
  PIN addrA1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 410.000 353.650 414.000 ;
    END
  END addrA1[5]
  PIN addrA1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 410.000 357.330 414.000 ;
    END
  END addrA1[6]
  PIN addrA1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 410.000 360.550 414.000 ;
    END
  END addrA1[7]
  PIN addrB0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END addrB0[0]
  PIN addrB0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 389.680 380.000 390.280 ;
    END
  END addrB0[1]
  PIN addrB0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 380.160 380.000 380.760 ;
    END
  END addrB0[2]
  PIN addrB0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 370.640 380.000 371.240 ;
    END
  END addrB0[3]
  PIN addrB0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 361.120 380.000 361.720 ;
    END
  END addrB0[4]
  PIN addrB0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 352.280 380.000 352.880 ;
    END
  END addrB0[5]
  PIN addrB0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 342.760 380.000 343.360 ;
    END
  END addrB0[6]
  PIN addrB0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 333.240 380.000 333.840 ;
    END
  END addrB0[7]
  PIN addrB0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 323.720 380.000 324.320 ;
    END
  END addrB0[8]
  PIN addrB1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 12.960 380.000 13.560 ;
    END
  END addrB1[0]
  PIN addrB1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 4.120 380.000 4.720 ;
    END
  END addrB1[1]
  PIN addrB1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END addrB1[2]
  PIN addrB1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END addrB1[3]
  PIN addrB1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 0.000 372.970 4.000 ;
    END
  END addrB1[4]
  PIN addrB1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END addrB1[5]
  PIN addrB1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END addrB1[6]
  PIN addrB1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END addrB1[7]
  PIN addrB1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END addrB1[8]
  PIN csbA0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END csbA0
  PIN csbA1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 410.000 378.030 414.000 ;
    END
  END csbA1
  PIN csbB0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 408.720 380.000 409.320 ;
    END
  END csbB0
  PIN csbB1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END csbB1
  PIN dinA0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 410.000 132.850 414.000 ;
    END
  END dinA0[0]
  PIN dinA0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 410.000 167.350 414.000 ;
    END
  END dinA0[10]
  PIN dinA0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 410.000 170.570 414.000 ;
    END
  END dinA0[11]
  PIN dinA0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 410.000 174.250 414.000 ;
    END
  END dinA0[12]
  PIN dinA0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 410.000 177.470 414.000 ;
    END
  END dinA0[13]
  PIN dinA0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 410.000 181.150 414.000 ;
    END
  END dinA0[14]
  PIN dinA0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 410.000 184.370 414.000 ;
    END
  END dinA0[15]
  PIN dinA0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 410.000 188.050 414.000 ;
    END
  END dinA0[16]
  PIN dinA0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 410.000 191.730 414.000 ;
    END
  END dinA0[17]
  PIN dinA0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 410.000 194.950 414.000 ;
    END
  END dinA0[18]
  PIN dinA0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 410.000 198.630 414.000 ;
    END
  END dinA0[19]
  PIN dinA0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 410.000 136.070 414.000 ;
    END
  END dinA0[1]
  PIN dinA0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 410.000 201.850 414.000 ;
    END
  END dinA0[20]
  PIN dinA0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 410.000 205.530 414.000 ;
    END
  END dinA0[21]
  PIN dinA0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 410.000 208.750 414.000 ;
    END
  END dinA0[22]
  PIN dinA0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 410.000 212.430 414.000 ;
    END
  END dinA0[23]
  PIN dinA0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 410.000 215.650 414.000 ;
    END
  END dinA0[24]
  PIN dinA0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 410.000 219.330 414.000 ;
    END
  END dinA0[25]
  PIN dinA0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 410.000 222.550 414.000 ;
    END
  END dinA0[26]
  PIN dinA0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 410.000 226.230 414.000 ;
    END
  END dinA0[27]
  PIN dinA0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 410.000 229.450 414.000 ;
    END
  END dinA0[28]
  PIN dinA0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 410.000 233.130 414.000 ;
    END
  END dinA0[29]
  PIN dinA0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 410.000 139.750 414.000 ;
    END
  END dinA0[2]
  PIN dinA0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 410.000 236.350 414.000 ;
    END
  END dinA0[30]
  PIN dinA0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 410.000 240.030 414.000 ;
    END
  END dinA0[31]
  PIN dinA0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 410.000 142.970 414.000 ;
    END
  END dinA0[3]
  PIN dinA0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 410.000 146.650 414.000 ;
    END
  END dinA0[4]
  PIN dinA0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 410.000 149.870 414.000 ;
    END
  END dinA0[5]
  PIN dinA0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 410.000 153.550 414.000 ;
    END
  END dinA0[6]
  PIN dinA0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 410.000 156.770 414.000 ;
    END
  END dinA0[7]
  PIN dinA0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 410.000 160.450 414.000 ;
    END
  END dinA0[8]
  PIN dinA0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 410.000 163.670 414.000 ;
    END
  END dinA0[9]
  PIN dinB0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END dinB0[0]
  PIN dinB0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END dinB0[10]
  PIN dinB0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END dinB0[11]
  PIN dinB0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END dinB0[12]
  PIN dinB0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END dinB0[13]
  PIN dinB0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END dinB0[14]
  PIN dinB0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END dinB0[15]
  PIN dinB0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END dinB0[16]
  PIN dinB0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END dinB0[17]
  PIN dinB0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END dinB0[18]
  PIN dinB0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END dinB0[19]
  PIN dinB0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END dinB0[1]
  PIN dinB0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END dinB0[20]
  PIN dinB0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END dinB0[21]
  PIN dinB0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END dinB0[22]
  PIN dinB0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END dinB0[23]
  PIN dinB0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END dinB0[24]
  PIN dinB0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END dinB0[25]
  PIN dinB0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END dinB0[26]
  PIN dinB0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END dinB0[27]
  PIN dinB0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END dinB0[28]
  PIN dinB0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END dinB0[29]
  PIN dinB0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END dinB0[2]
  PIN dinB0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END dinB0[30]
  PIN dinB0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END dinB0[31]
  PIN dinB0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END dinB0[3]
  PIN dinB0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END dinB0[4]
  PIN dinB0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END dinB0[5]
  PIN dinB0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END dinB0[6]
  PIN dinB0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END dinB0[7]
  PIN dinB0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END dinB0[8]
  PIN dinB0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END dinB0[9]
  PIN sram12_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END sram12_dout0[0]
  PIN sram12_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END sram12_dout0[10]
  PIN sram12_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END sram12_dout0[11]
  PIN sram12_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END sram12_dout0[12]
  PIN sram12_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END sram12_dout0[13]
  PIN sram12_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END sram12_dout0[14]
  PIN sram12_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END sram12_dout0[15]
  PIN sram12_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END sram12_dout0[16]
  PIN sram12_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END sram12_dout0[17]
  PIN sram12_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END sram12_dout0[18]
  PIN sram12_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END sram12_dout0[19]
  PIN sram12_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END sram12_dout0[1]
  PIN sram12_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END sram12_dout0[20]
  PIN sram12_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END sram12_dout0[21]
  PIN sram12_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END sram12_dout0[22]
  PIN sram12_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END sram12_dout0[23]
  PIN sram12_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END sram12_dout0[24]
  PIN sram12_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END sram12_dout0[25]
  PIN sram12_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END sram12_dout0[26]
  PIN sram12_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END sram12_dout0[27]
  PIN sram12_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END sram12_dout0[28]
  PIN sram12_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END sram12_dout0[29]
  PIN sram12_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END sram12_dout0[2]
  PIN sram12_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END sram12_dout0[30]
  PIN sram12_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END sram12_dout0[31]
  PIN sram12_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END sram12_dout0[3]
  PIN sram12_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END sram12_dout0[4]
  PIN sram12_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END sram12_dout0[5]
  PIN sram12_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END sram12_dout0[6]
  PIN sram12_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END sram12_dout0[7]
  PIN sram12_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END sram12_dout0[8]
  PIN sram12_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END sram12_dout0[9]
  PIN sram12_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 22.480 380.000 23.080 ;
    END
  END sram12_dout1[0]
  PIN sram12_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 117.000 380.000 117.600 ;
    END
  END sram12_dout1[10]
  PIN sram12_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 125.840 380.000 126.440 ;
    END
  END sram12_dout1[11]
  PIN sram12_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 135.360 380.000 135.960 ;
    END
  END sram12_dout1[12]
  PIN sram12_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 144.880 380.000 145.480 ;
    END
  END sram12_dout1[13]
  PIN sram12_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 154.400 380.000 155.000 ;
    END
  END sram12_dout1[14]
  PIN sram12_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 163.920 380.000 164.520 ;
    END
  END sram12_dout1[15]
  PIN sram12_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 173.440 380.000 174.040 ;
    END
  END sram12_dout1[16]
  PIN sram12_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 182.280 380.000 182.880 ;
    END
  END sram12_dout1[17]
  PIN sram12_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 191.800 380.000 192.400 ;
    END
  END sram12_dout1[18]
  PIN sram12_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 201.320 380.000 201.920 ;
    END
  END sram12_dout1[19]
  PIN sram12_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 32.000 380.000 32.600 ;
    END
  END sram12_dout1[1]
  PIN sram12_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 210.840 380.000 211.440 ;
    END
  END sram12_dout1[20]
  PIN sram12_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 220.360 380.000 220.960 ;
    END
  END sram12_dout1[21]
  PIN sram12_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 229.880 380.000 230.480 ;
    END
  END sram12_dout1[22]
  PIN sram12_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 239.400 380.000 240.000 ;
    END
  END sram12_dout1[23]
  PIN sram12_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 248.240 380.000 248.840 ;
    END
  END sram12_dout1[24]
  PIN sram12_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 257.760 380.000 258.360 ;
    END
  END sram12_dout1[25]
  PIN sram12_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 267.280 380.000 267.880 ;
    END
  END sram12_dout1[26]
  PIN sram12_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 276.800 380.000 277.400 ;
    END
  END sram12_dout1[27]
  PIN sram12_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 286.320 380.000 286.920 ;
    END
  END sram12_dout1[28]
  PIN sram12_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 295.840 380.000 296.440 ;
    END
  END sram12_dout1[29]
  PIN sram12_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 41.520 380.000 42.120 ;
    END
  END sram12_dout1[2]
  PIN sram12_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 304.680 380.000 305.280 ;
    END
  END sram12_dout1[30]
  PIN sram12_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 314.200 380.000 314.800 ;
    END
  END sram12_dout1[31]
  PIN sram12_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 51.040 380.000 51.640 ;
    END
  END sram12_dout1[3]
  PIN sram12_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 60.560 380.000 61.160 ;
    END
  END sram12_dout1[4]
  PIN sram12_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 69.400 380.000 70.000 ;
    END
  END sram12_dout1[5]
  PIN sram12_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 78.920 380.000 79.520 ;
    END
  END sram12_dout1[6]
  PIN sram12_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 88.440 380.000 89.040 ;
    END
  END sram12_dout1[7]
  PIN sram12_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 97.960 380.000 98.560 ;
    END
  END sram12_dout1[8]
  PIN sram12_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 107.480 380.000 108.080 ;
    END
  END sram12_dout1[9]
  PIN sram1_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 410.000 243.250 414.000 ;
    END
  END sram1_dout0[0]
  PIN sram1_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 410.000 277.750 414.000 ;
    END
  END sram1_dout0[10]
  PIN sram1_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 410.000 281.430 414.000 ;
    END
  END sram1_dout0[11]
  PIN sram1_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 410.000 284.650 414.000 ;
    END
  END sram1_dout0[12]
  PIN sram1_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 410.000 288.330 414.000 ;
    END
  END sram1_dout0[13]
  PIN sram1_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 410.000 291.550 414.000 ;
    END
  END sram1_dout0[14]
  PIN sram1_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 410.000 295.230 414.000 ;
    END
  END sram1_dout0[15]
  PIN sram1_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 410.000 298.450 414.000 ;
    END
  END sram1_dout0[16]
  PIN sram1_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 410.000 302.130 414.000 ;
    END
  END sram1_dout0[17]
  PIN sram1_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 410.000 305.350 414.000 ;
    END
  END sram1_dout0[18]
  PIN sram1_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 410.000 309.030 414.000 ;
    END
  END sram1_dout0[19]
  PIN sram1_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 410.000 246.930 414.000 ;
    END
  END sram1_dout0[1]
  PIN sram1_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 410.000 312.250 414.000 ;
    END
  END sram1_dout0[20]
  PIN sram1_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 410.000 315.930 414.000 ;
    END
  END sram1_dout0[21]
  PIN sram1_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 410.000 319.150 414.000 ;
    END
  END sram1_dout0[22]
  PIN sram1_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 410.000 322.830 414.000 ;
    END
  END sram1_dout0[23]
  PIN sram1_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 410.000 326.050 414.000 ;
    END
  END sram1_dout0[24]
  PIN sram1_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 410.000 329.730 414.000 ;
    END
  END sram1_dout0[25]
  PIN sram1_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 410.000 332.950 414.000 ;
    END
  END sram1_dout0[26]
  PIN sram1_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 410.000 336.630 414.000 ;
    END
  END sram1_dout0[27]
  PIN sram1_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 410.000 339.850 414.000 ;
    END
  END sram1_dout0[28]
  PIN sram1_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 410.000 343.530 414.000 ;
    END
  END sram1_dout0[29]
  PIN sram1_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 410.000 250.150 414.000 ;
    END
  END sram1_dout0[2]
  PIN sram1_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 410.000 346.750 414.000 ;
    END
  END sram1_dout0[30]
  PIN sram1_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 410.000 350.430 414.000 ;
    END
  END sram1_dout0[31]
  PIN sram1_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 410.000 253.830 414.000 ;
    END
  END sram1_dout0[3]
  PIN sram1_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 410.000 257.050 414.000 ;
    END
  END sram1_dout0[4]
  PIN sram1_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 410.000 260.730 414.000 ;
    END
  END sram1_dout0[5]
  PIN sram1_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 410.000 263.950 414.000 ;
    END
  END sram1_dout0[6]
  PIN sram1_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 410.000 267.630 414.000 ;
    END
  END sram1_dout0[7]
  PIN sram1_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 410.000 270.850 414.000 ;
    END
  END sram1_dout0[8]
  PIN sram1_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 410.000 274.530 414.000 ;
    END
  END sram1_dout0[9]
  PIN sram1_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 410.000 1.750 414.000 ;
    END
  END sram1_dout1[0]
  PIN sram1_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 410.000 36.250 414.000 ;
    END
  END sram1_dout1[10]
  PIN sram1_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 410.000 39.470 414.000 ;
    END
  END sram1_dout1[11]
  PIN sram1_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 410.000 43.150 414.000 ;
    END
  END sram1_dout1[12]
  PIN sram1_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 410.000 46.370 414.000 ;
    END
  END sram1_dout1[13]
  PIN sram1_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 410.000 50.050 414.000 ;
    END
  END sram1_dout1[14]
  PIN sram1_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 410.000 53.270 414.000 ;
    END
  END sram1_dout1[15]
  PIN sram1_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 410.000 56.950 414.000 ;
    END
  END sram1_dout1[16]
  PIN sram1_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 410.000 60.170 414.000 ;
    END
  END sram1_dout1[17]
  PIN sram1_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 410.000 63.850 414.000 ;
    END
  END sram1_dout1[18]
  PIN sram1_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 410.000 67.070 414.000 ;
    END
  END sram1_dout1[19]
  PIN sram1_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 410.000 4.970 414.000 ;
    END
  END sram1_dout1[1]
  PIN sram1_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 410.000 70.750 414.000 ;
    END
  END sram1_dout1[20]
  PIN sram1_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 410.000 73.970 414.000 ;
    END
  END sram1_dout1[21]
  PIN sram1_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 410.000 77.650 414.000 ;
    END
  END sram1_dout1[22]
  PIN sram1_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 410.000 80.870 414.000 ;
    END
  END sram1_dout1[23]
  PIN sram1_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 410.000 84.550 414.000 ;
    END
  END sram1_dout1[24]
  PIN sram1_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 410.000 87.770 414.000 ;
    END
  END sram1_dout1[25]
  PIN sram1_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 410.000 91.450 414.000 ;
    END
  END sram1_dout1[26]
  PIN sram1_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 410.000 94.670 414.000 ;
    END
  END sram1_dout1[27]
  PIN sram1_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 410.000 98.350 414.000 ;
    END
  END sram1_dout1[28]
  PIN sram1_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 410.000 101.570 414.000 ;
    END
  END sram1_dout1[29]
  PIN sram1_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 410.000 8.650 414.000 ;
    END
  END sram1_dout1[2]
  PIN sram1_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 410.000 105.250 414.000 ;
    END
  END sram1_dout1[30]
  PIN sram1_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 410.000 108.470 414.000 ;
    END
  END sram1_dout1[31]
  PIN sram1_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 410.000 11.870 414.000 ;
    END
  END sram1_dout1[3]
  PIN sram1_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 410.000 15.550 414.000 ;
    END
  END sram1_dout1[4]
  PIN sram1_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 410.000 18.770 414.000 ;
    END
  END sram1_dout1[5]
  PIN sram1_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 410.000 22.450 414.000 ;
    END
  END sram1_dout1[6]
  PIN sram1_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 410.000 25.670 414.000 ;
    END
  END sram1_dout1[7]
  PIN sram1_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 410.000 29.350 414.000 ;
    END
  END sram1_dout1[8]
  PIN sram1_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 410.000 32.570 414.000 ;
    END
  END sram1_dout1[9]
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 402.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 402.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 402.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 402.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 402.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END wbs_we_i
  PIN webA
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END webA
  PIN webB
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.000 399.200 380.000 399.800 ;
    END
  END webB
  PIN wmaskA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 410.000 119.050 414.000 ;
    END
  END wmaskA[0]
  PIN wmaskA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 410.000 122.270 414.000 ;
    END
  END wmaskA[1]
  PIN wmaskA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 410.000 125.950 414.000 ;
    END
  END wmaskA[2]
  PIN wmaskA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 410.000 129.170 414.000 ;
    END
  END wmaskA[3]
  PIN wmaskB[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END wmaskB[0]
  PIN wmaskB[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END wmaskB[1]
  PIN wmaskB[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END wmaskB[2]
  PIN wmaskB[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END wmaskB[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 374.440 402.645 ;
      LAYER met1 ;
        RECT 0.070 0.040 379.890 405.240 ;
      LAYER met2 ;
        RECT 0.100 409.720 1.190 410.450 ;
        RECT 2.030 409.720 4.410 410.450 ;
        RECT 5.250 409.720 8.090 410.450 ;
        RECT 8.930 409.720 11.310 410.450 ;
        RECT 12.150 409.720 14.990 410.450 ;
        RECT 15.830 409.720 18.210 410.450 ;
        RECT 19.050 409.720 21.890 410.450 ;
        RECT 22.730 409.720 25.110 410.450 ;
        RECT 25.950 409.720 28.790 410.450 ;
        RECT 29.630 409.720 32.010 410.450 ;
        RECT 32.850 409.720 35.690 410.450 ;
        RECT 36.530 409.720 38.910 410.450 ;
        RECT 39.750 409.720 42.590 410.450 ;
        RECT 43.430 409.720 45.810 410.450 ;
        RECT 46.650 409.720 49.490 410.450 ;
        RECT 50.330 409.720 52.710 410.450 ;
        RECT 53.550 409.720 56.390 410.450 ;
        RECT 57.230 409.720 59.610 410.450 ;
        RECT 60.450 409.720 63.290 410.450 ;
        RECT 64.130 409.720 66.510 410.450 ;
        RECT 67.350 409.720 70.190 410.450 ;
        RECT 71.030 409.720 73.410 410.450 ;
        RECT 74.250 409.720 77.090 410.450 ;
        RECT 77.930 409.720 80.310 410.450 ;
        RECT 81.150 409.720 83.990 410.450 ;
        RECT 84.830 409.720 87.210 410.450 ;
        RECT 88.050 409.720 90.890 410.450 ;
        RECT 91.730 409.720 94.110 410.450 ;
        RECT 94.950 409.720 97.790 410.450 ;
        RECT 98.630 409.720 101.010 410.450 ;
        RECT 101.850 409.720 104.690 410.450 ;
        RECT 105.530 409.720 107.910 410.450 ;
        RECT 108.750 409.720 111.590 410.450 ;
        RECT 112.430 409.720 114.810 410.450 ;
        RECT 115.650 409.720 118.490 410.450 ;
        RECT 119.330 409.720 121.710 410.450 ;
        RECT 122.550 409.720 125.390 410.450 ;
        RECT 126.230 409.720 128.610 410.450 ;
        RECT 129.450 409.720 132.290 410.450 ;
        RECT 133.130 409.720 135.510 410.450 ;
        RECT 136.350 409.720 139.190 410.450 ;
        RECT 140.030 409.720 142.410 410.450 ;
        RECT 143.250 409.720 146.090 410.450 ;
        RECT 146.930 409.720 149.310 410.450 ;
        RECT 150.150 409.720 152.990 410.450 ;
        RECT 153.830 409.720 156.210 410.450 ;
        RECT 157.050 409.720 159.890 410.450 ;
        RECT 160.730 409.720 163.110 410.450 ;
        RECT 163.950 409.720 166.790 410.450 ;
        RECT 167.630 409.720 170.010 410.450 ;
        RECT 170.850 409.720 173.690 410.450 ;
        RECT 174.530 409.720 176.910 410.450 ;
        RECT 177.750 409.720 180.590 410.450 ;
        RECT 181.430 409.720 183.810 410.450 ;
        RECT 184.650 409.720 187.490 410.450 ;
        RECT 188.330 409.720 191.170 410.450 ;
        RECT 192.010 409.720 194.390 410.450 ;
        RECT 195.230 409.720 198.070 410.450 ;
        RECT 198.910 409.720 201.290 410.450 ;
        RECT 202.130 409.720 204.970 410.450 ;
        RECT 205.810 409.720 208.190 410.450 ;
        RECT 209.030 409.720 211.870 410.450 ;
        RECT 212.710 409.720 215.090 410.450 ;
        RECT 215.930 409.720 218.770 410.450 ;
        RECT 219.610 409.720 221.990 410.450 ;
        RECT 222.830 409.720 225.670 410.450 ;
        RECT 226.510 409.720 228.890 410.450 ;
        RECT 229.730 409.720 232.570 410.450 ;
        RECT 233.410 409.720 235.790 410.450 ;
        RECT 236.630 409.720 239.470 410.450 ;
        RECT 240.310 409.720 242.690 410.450 ;
        RECT 243.530 409.720 246.370 410.450 ;
        RECT 247.210 409.720 249.590 410.450 ;
        RECT 250.430 409.720 253.270 410.450 ;
        RECT 254.110 409.720 256.490 410.450 ;
        RECT 257.330 409.720 260.170 410.450 ;
        RECT 261.010 409.720 263.390 410.450 ;
        RECT 264.230 409.720 267.070 410.450 ;
        RECT 267.910 409.720 270.290 410.450 ;
        RECT 271.130 409.720 273.970 410.450 ;
        RECT 274.810 409.720 277.190 410.450 ;
        RECT 278.030 409.720 280.870 410.450 ;
        RECT 281.710 409.720 284.090 410.450 ;
        RECT 284.930 409.720 287.770 410.450 ;
        RECT 288.610 409.720 290.990 410.450 ;
        RECT 291.830 409.720 294.670 410.450 ;
        RECT 295.510 409.720 297.890 410.450 ;
        RECT 298.730 409.720 301.570 410.450 ;
        RECT 302.410 409.720 304.790 410.450 ;
        RECT 305.630 409.720 308.470 410.450 ;
        RECT 309.310 409.720 311.690 410.450 ;
        RECT 312.530 409.720 315.370 410.450 ;
        RECT 316.210 409.720 318.590 410.450 ;
        RECT 319.430 409.720 322.270 410.450 ;
        RECT 323.110 409.720 325.490 410.450 ;
        RECT 326.330 409.720 329.170 410.450 ;
        RECT 330.010 409.720 332.390 410.450 ;
        RECT 333.230 409.720 336.070 410.450 ;
        RECT 336.910 409.720 339.290 410.450 ;
        RECT 340.130 409.720 342.970 410.450 ;
        RECT 343.810 409.720 346.190 410.450 ;
        RECT 347.030 409.720 349.870 410.450 ;
        RECT 350.710 409.720 353.090 410.450 ;
        RECT 353.930 409.720 356.770 410.450 ;
        RECT 357.610 409.720 359.990 410.450 ;
        RECT 360.830 409.720 363.670 410.450 ;
        RECT 364.510 409.720 366.890 410.450 ;
        RECT 367.730 409.720 370.570 410.450 ;
        RECT 371.410 409.720 373.790 410.450 ;
        RECT 374.630 409.720 377.470 410.450 ;
        RECT 378.310 409.720 379.870 410.450 ;
        RECT 0.100 4.280 379.870 409.720 ;
        RECT 0.100 0.010 0.730 4.280 ;
        RECT 1.570 0.010 2.570 4.280 ;
        RECT 3.410 0.010 4.410 4.280 ;
        RECT 5.250 0.010 6.710 4.280 ;
        RECT 7.550 0.010 8.550 4.280 ;
        RECT 9.390 0.010 10.850 4.280 ;
        RECT 11.690 0.010 12.690 4.280 ;
        RECT 13.530 0.010 14.990 4.280 ;
        RECT 15.830 0.010 16.830 4.280 ;
        RECT 17.670 0.010 18.670 4.280 ;
        RECT 19.510 0.010 20.970 4.280 ;
        RECT 21.810 0.010 22.810 4.280 ;
        RECT 23.650 0.010 25.110 4.280 ;
        RECT 25.950 0.010 26.950 4.280 ;
        RECT 27.790 0.010 29.250 4.280 ;
        RECT 30.090 0.010 31.090 4.280 ;
        RECT 31.930 0.010 33.390 4.280 ;
        RECT 34.230 0.010 35.230 4.280 ;
        RECT 36.070 0.010 37.070 4.280 ;
        RECT 37.910 0.010 39.370 4.280 ;
        RECT 40.210 0.010 41.210 4.280 ;
        RECT 42.050 0.010 43.510 4.280 ;
        RECT 44.350 0.010 45.350 4.280 ;
        RECT 46.190 0.010 47.650 4.280 ;
        RECT 48.490 0.010 49.490 4.280 ;
        RECT 50.330 0.010 51.790 4.280 ;
        RECT 52.630 0.010 53.630 4.280 ;
        RECT 54.470 0.010 55.470 4.280 ;
        RECT 56.310 0.010 57.770 4.280 ;
        RECT 58.610 0.010 59.610 4.280 ;
        RECT 60.450 0.010 61.910 4.280 ;
        RECT 62.750 0.010 63.750 4.280 ;
        RECT 64.590 0.010 66.050 4.280 ;
        RECT 66.890 0.010 67.890 4.280 ;
        RECT 68.730 0.010 69.730 4.280 ;
        RECT 70.570 0.010 72.030 4.280 ;
        RECT 72.870 0.010 73.870 4.280 ;
        RECT 74.710 0.010 76.170 4.280 ;
        RECT 77.010 0.010 78.010 4.280 ;
        RECT 78.850 0.010 80.310 4.280 ;
        RECT 81.150 0.010 82.150 4.280 ;
        RECT 82.990 0.010 84.450 4.280 ;
        RECT 85.290 0.010 86.290 4.280 ;
        RECT 87.130 0.010 88.130 4.280 ;
        RECT 88.970 0.010 90.430 4.280 ;
        RECT 91.270 0.010 92.270 4.280 ;
        RECT 93.110 0.010 94.570 4.280 ;
        RECT 95.410 0.010 96.410 4.280 ;
        RECT 97.250 0.010 98.710 4.280 ;
        RECT 99.550 0.010 100.550 4.280 ;
        RECT 101.390 0.010 102.850 4.280 ;
        RECT 103.690 0.010 104.690 4.280 ;
        RECT 105.530 0.010 106.530 4.280 ;
        RECT 107.370 0.010 108.830 4.280 ;
        RECT 109.670 0.010 110.670 4.280 ;
        RECT 111.510 0.010 112.970 4.280 ;
        RECT 113.810 0.010 114.810 4.280 ;
        RECT 115.650 0.010 117.110 4.280 ;
        RECT 117.950 0.010 118.950 4.280 ;
        RECT 119.790 0.010 121.250 4.280 ;
        RECT 122.090 0.010 123.090 4.280 ;
        RECT 123.930 0.010 124.930 4.280 ;
        RECT 125.770 0.010 127.230 4.280 ;
        RECT 128.070 0.010 129.070 4.280 ;
        RECT 129.910 0.010 131.370 4.280 ;
        RECT 132.210 0.010 133.210 4.280 ;
        RECT 134.050 0.010 135.510 4.280 ;
        RECT 136.350 0.010 137.350 4.280 ;
        RECT 138.190 0.010 139.190 4.280 ;
        RECT 140.030 0.010 141.490 4.280 ;
        RECT 142.330 0.010 143.330 4.280 ;
        RECT 144.170 0.010 145.630 4.280 ;
        RECT 146.470 0.010 147.470 4.280 ;
        RECT 148.310 0.010 149.770 4.280 ;
        RECT 150.610 0.010 151.610 4.280 ;
        RECT 152.450 0.010 153.910 4.280 ;
        RECT 154.750 0.010 155.750 4.280 ;
        RECT 156.590 0.010 157.590 4.280 ;
        RECT 158.430 0.010 159.890 4.280 ;
        RECT 160.730 0.010 161.730 4.280 ;
        RECT 162.570 0.010 164.030 4.280 ;
        RECT 164.870 0.010 165.870 4.280 ;
        RECT 166.710 0.010 168.170 4.280 ;
        RECT 169.010 0.010 170.010 4.280 ;
        RECT 170.850 0.010 172.310 4.280 ;
        RECT 173.150 0.010 174.150 4.280 ;
        RECT 174.990 0.010 175.990 4.280 ;
        RECT 176.830 0.010 178.290 4.280 ;
        RECT 179.130 0.010 180.130 4.280 ;
        RECT 180.970 0.010 182.430 4.280 ;
        RECT 183.270 0.010 184.270 4.280 ;
        RECT 185.110 0.010 186.570 4.280 ;
        RECT 187.410 0.010 188.410 4.280 ;
        RECT 189.250 0.010 190.710 4.280 ;
        RECT 191.550 0.010 192.550 4.280 ;
        RECT 193.390 0.010 194.390 4.280 ;
        RECT 195.230 0.010 196.690 4.280 ;
        RECT 197.530 0.010 198.530 4.280 ;
        RECT 199.370 0.010 200.830 4.280 ;
        RECT 201.670 0.010 202.670 4.280 ;
        RECT 203.510 0.010 204.970 4.280 ;
        RECT 205.810 0.010 206.810 4.280 ;
        RECT 207.650 0.010 208.650 4.280 ;
        RECT 209.490 0.010 210.950 4.280 ;
        RECT 211.790 0.010 212.790 4.280 ;
        RECT 213.630 0.010 215.090 4.280 ;
        RECT 215.930 0.010 216.930 4.280 ;
        RECT 217.770 0.010 219.230 4.280 ;
        RECT 220.070 0.010 221.070 4.280 ;
        RECT 221.910 0.010 223.370 4.280 ;
        RECT 224.210 0.010 225.210 4.280 ;
        RECT 226.050 0.010 227.050 4.280 ;
        RECT 227.890 0.010 229.350 4.280 ;
        RECT 230.190 0.010 231.190 4.280 ;
        RECT 232.030 0.010 233.490 4.280 ;
        RECT 234.330 0.010 235.330 4.280 ;
        RECT 236.170 0.010 237.630 4.280 ;
        RECT 238.470 0.010 239.470 4.280 ;
        RECT 240.310 0.010 241.770 4.280 ;
        RECT 242.610 0.010 243.610 4.280 ;
        RECT 244.450 0.010 245.450 4.280 ;
        RECT 246.290 0.010 247.750 4.280 ;
        RECT 248.590 0.010 249.590 4.280 ;
        RECT 250.430 0.010 251.890 4.280 ;
        RECT 252.730 0.010 253.730 4.280 ;
        RECT 254.570 0.010 256.030 4.280 ;
        RECT 256.870 0.010 257.870 4.280 ;
        RECT 258.710 0.010 259.710 4.280 ;
        RECT 260.550 0.010 262.010 4.280 ;
        RECT 262.850 0.010 263.850 4.280 ;
        RECT 264.690 0.010 266.150 4.280 ;
        RECT 266.990 0.010 267.990 4.280 ;
        RECT 268.830 0.010 270.290 4.280 ;
        RECT 271.130 0.010 272.130 4.280 ;
        RECT 272.970 0.010 274.430 4.280 ;
        RECT 275.270 0.010 276.270 4.280 ;
        RECT 277.110 0.010 278.110 4.280 ;
        RECT 278.950 0.010 280.410 4.280 ;
        RECT 281.250 0.010 282.250 4.280 ;
        RECT 283.090 0.010 284.550 4.280 ;
        RECT 285.390 0.010 286.390 4.280 ;
        RECT 287.230 0.010 288.690 4.280 ;
        RECT 289.530 0.010 290.530 4.280 ;
        RECT 291.370 0.010 292.830 4.280 ;
        RECT 293.670 0.010 294.670 4.280 ;
        RECT 295.510 0.010 296.510 4.280 ;
        RECT 297.350 0.010 298.810 4.280 ;
        RECT 299.650 0.010 300.650 4.280 ;
        RECT 301.490 0.010 302.950 4.280 ;
        RECT 303.790 0.010 304.790 4.280 ;
        RECT 305.630 0.010 307.090 4.280 ;
        RECT 307.930 0.010 308.930 4.280 ;
        RECT 309.770 0.010 311.230 4.280 ;
        RECT 312.070 0.010 313.070 4.280 ;
        RECT 313.910 0.010 314.910 4.280 ;
        RECT 315.750 0.010 317.210 4.280 ;
        RECT 318.050 0.010 319.050 4.280 ;
        RECT 319.890 0.010 321.350 4.280 ;
        RECT 322.190 0.010 323.190 4.280 ;
        RECT 324.030 0.010 325.490 4.280 ;
        RECT 326.330 0.010 327.330 4.280 ;
        RECT 328.170 0.010 329.170 4.280 ;
        RECT 330.010 0.010 331.470 4.280 ;
        RECT 332.310 0.010 333.310 4.280 ;
        RECT 334.150 0.010 335.610 4.280 ;
        RECT 336.450 0.010 337.450 4.280 ;
        RECT 338.290 0.010 339.750 4.280 ;
        RECT 340.590 0.010 341.590 4.280 ;
        RECT 342.430 0.010 343.890 4.280 ;
        RECT 344.730 0.010 345.730 4.280 ;
        RECT 346.570 0.010 347.570 4.280 ;
        RECT 348.410 0.010 349.870 4.280 ;
        RECT 350.710 0.010 351.710 4.280 ;
        RECT 352.550 0.010 354.010 4.280 ;
        RECT 354.850 0.010 355.850 4.280 ;
        RECT 356.690 0.010 358.150 4.280 ;
        RECT 358.990 0.010 359.990 4.280 ;
        RECT 360.830 0.010 362.290 4.280 ;
        RECT 363.130 0.010 364.130 4.280 ;
        RECT 364.970 0.010 365.970 4.280 ;
        RECT 366.810 0.010 368.270 4.280 ;
        RECT 369.110 0.010 370.110 4.280 ;
        RECT 370.950 0.010 372.410 4.280 ;
        RECT 373.250 0.010 374.250 4.280 ;
        RECT 375.090 0.010 376.550 4.280 ;
        RECT 377.390 0.010 378.390 4.280 ;
        RECT 379.230 0.010 379.870 4.280 ;
      LAYER met3 ;
        RECT 4.000 408.320 375.600 409.185 ;
        RECT 4.000 400.200 379.895 408.320 ;
        RECT 4.000 398.800 375.600 400.200 ;
        RECT 4.000 391.360 379.895 398.800 ;
        RECT 4.400 390.680 379.895 391.360 ;
        RECT 4.400 389.960 375.600 390.680 ;
        RECT 4.000 389.280 375.600 389.960 ;
        RECT 4.000 381.160 379.895 389.280 ;
        RECT 4.000 379.760 375.600 381.160 ;
        RECT 4.000 371.640 379.895 379.760 ;
        RECT 4.000 370.240 375.600 371.640 ;
        RECT 4.000 362.120 379.895 370.240 ;
        RECT 4.000 360.720 375.600 362.120 ;
        RECT 4.000 353.280 379.895 360.720 ;
        RECT 4.000 351.880 375.600 353.280 ;
        RECT 4.000 345.120 379.895 351.880 ;
        RECT 4.400 343.760 379.895 345.120 ;
        RECT 4.400 343.720 375.600 343.760 ;
        RECT 4.000 342.360 375.600 343.720 ;
        RECT 4.000 334.240 379.895 342.360 ;
        RECT 4.000 332.840 375.600 334.240 ;
        RECT 4.000 324.720 379.895 332.840 ;
        RECT 4.000 323.320 375.600 324.720 ;
        RECT 4.000 315.200 379.895 323.320 ;
        RECT 4.000 313.800 375.600 315.200 ;
        RECT 4.000 305.680 379.895 313.800 ;
        RECT 4.000 304.280 375.600 305.680 ;
        RECT 4.000 299.560 379.895 304.280 ;
        RECT 4.400 298.160 379.895 299.560 ;
        RECT 4.000 296.840 379.895 298.160 ;
        RECT 4.000 295.440 375.600 296.840 ;
        RECT 4.000 287.320 379.895 295.440 ;
        RECT 4.000 285.920 375.600 287.320 ;
        RECT 4.000 277.800 379.895 285.920 ;
        RECT 4.000 276.400 375.600 277.800 ;
        RECT 4.000 268.280 379.895 276.400 ;
        RECT 4.000 266.880 375.600 268.280 ;
        RECT 4.000 258.760 379.895 266.880 ;
        RECT 4.000 257.360 375.600 258.760 ;
        RECT 4.000 253.320 379.895 257.360 ;
        RECT 4.400 251.920 379.895 253.320 ;
        RECT 4.000 249.240 379.895 251.920 ;
        RECT 4.000 247.840 375.600 249.240 ;
        RECT 4.000 240.400 379.895 247.840 ;
        RECT 4.000 239.000 375.600 240.400 ;
        RECT 4.000 230.880 379.895 239.000 ;
        RECT 4.000 229.480 375.600 230.880 ;
        RECT 4.000 221.360 379.895 229.480 ;
        RECT 4.000 219.960 375.600 221.360 ;
        RECT 4.000 211.840 379.895 219.960 ;
        RECT 4.000 210.440 375.600 211.840 ;
        RECT 4.000 207.080 379.895 210.440 ;
        RECT 4.400 205.680 379.895 207.080 ;
        RECT 4.000 202.320 379.895 205.680 ;
        RECT 4.000 200.920 375.600 202.320 ;
        RECT 4.000 192.800 379.895 200.920 ;
        RECT 4.000 191.400 375.600 192.800 ;
        RECT 4.000 183.280 379.895 191.400 ;
        RECT 4.000 181.880 375.600 183.280 ;
        RECT 4.000 174.440 379.895 181.880 ;
        RECT 4.000 173.040 375.600 174.440 ;
        RECT 4.000 164.920 379.895 173.040 ;
        RECT 4.000 163.520 375.600 164.920 ;
        RECT 4.000 161.520 379.895 163.520 ;
        RECT 4.400 160.120 379.895 161.520 ;
        RECT 4.000 155.400 379.895 160.120 ;
        RECT 4.000 154.000 375.600 155.400 ;
        RECT 4.000 145.880 379.895 154.000 ;
        RECT 4.000 144.480 375.600 145.880 ;
        RECT 4.000 136.360 379.895 144.480 ;
        RECT 4.000 134.960 375.600 136.360 ;
        RECT 4.000 126.840 379.895 134.960 ;
        RECT 4.000 125.440 375.600 126.840 ;
        RECT 4.000 118.000 379.895 125.440 ;
        RECT 4.000 116.600 375.600 118.000 ;
        RECT 4.000 115.280 379.895 116.600 ;
        RECT 4.400 113.880 379.895 115.280 ;
        RECT 4.000 108.480 379.895 113.880 ;
        RECT 4.000 107.080 375.600 108.480 ;
        RECT 4.000 98.960 379.895 107.080 ;
        RECT 4.000 97.560 375.600 98.960 ;
        RECT 4.000 89.440 379.895 97.560 ;
        RECT 4.000 88.040 375.600 89.440 ;
        RECT 4.000 79.920 379.895 88.040 ;
        RECT 4.000 78.520 375.600 79.920 ;
        RECT 4.000 70.400 379.895 78.520 ;
        RECT 4.000 69.040 375.600 70.400 ;
        RECT 4.400 69.000 375.600 69.040 ;
        RECT 4.400 67.640 379.895 69.000 ;
        RECT 4.000 61.560 379.895 67.640 ;
        RECT 4.000 60.160 375.600 61.560 ;
        RECT 4.000 52.040 379.895 60.160 ;
        RECT 4.000 50.640 375.600 52.040 ;
        RECT 4.000 42.520 379.895 50.640 ;
        RECT 4.000 41.120 375.600 42.520 ;
        RECT 4.000 33.000 379.895 41.120 ;
        RECT 4.000 31.600 375.600 33.000 ;
        RECT 4.000 23.480 379.895 31.600 ;
        RECT 4.400 22.080 375.600 23.480 ;
        RECT 4.000 13.960 379.895 22.080 ;
        RECT 4.000 12.560 375.600 13.960 ;
        RECT 4.000 5.120 379.895 12.560 ;
        RECT 4.000 3.720 375.600 5.120 ;
        RECT 4.000 0.175 379.895 3.720 ;
      LAYER met4 ;
        RECT 8.575 403.200 379.665 403.745 ;
        RECT 8.575 10.240 20.640 403.200 ;
        RECT 23.040 10.240 97.440 403.200 ;
        RECT 99.840 10.240 174.240 403.200 ;
        RECT 176.640 10.240 251.040 403.200 ;
        RECT 253.440 10.240 327.840 403.200 ;
        RECT 330.240 10.240 379.665 403.200 ;
        RECT 8.575 0.175 379.665 10.240 ;
  END
END user_project
END LIBRARY

