magic
tech sky130A
magscale 1 2
timestamp 1647358929
<< obsli1 >>
rect 20704 16159 94488 94529
<< obsm1 >>
rect 1670 8 582438 189236
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 110 536 583432 189242
rect 110 2 486 536
rect 710 2 1590 536
rect 1814 2 2786 536
rect 3010 2 3982 536
rect 4206 2 5178 536
rect 5402 2 6374 536
rect 6598 2 7570 536
rect 7794 2 8674 536
rect 8898 2 9870 536
rect 10094 2 11066 536
rect 11290 2 12262 536
rect 12486 2 13458 536
rect 13682 2 14654 536
rect 14878 2 15850 536
rect 16074 2 16954 536
rect 17178 2 18150 536
rect 18374 2 19346 536
rect 19570 2 20542 536
rect 20766 2 21738 536
rect 21962 2 22934 536
rect 23158 2 24130 536
rect 24354 2 25234 536
rect 25458 2 26430 536
rect 26654 2 27626 536
rect 27850 2 28822 536
rect 29046 2 30018 536
rect 30242 2 31214 536
rect 31438 2 32318 536
rect 32542 2 33514 536
rect 33738 2 34710 536
rect 34934 2 35906 536
rect 36130 2 37102 536
rect 37326 2 38298 536
rect 38522 2 39494 536
rect 39718 2 40598 536
rect 40822 2 41794 536
rect 42018 2 42990 536
rect 43214 2 44186 536
rect 44410 2 45382 536
rect 45606 2 46578 536
rect 46802 2 47774 536
rect 47998 2 48878 536
rect 49102 2 50074 536
rect 50298 2 51270 536
rect 51494 2 52466 536
rect 52690 2 53662 536
rect 53886 2 54858 536
rect 55082 2 55962 536
rect 56186 2 57158 536
rect 57382 2 58354 536
rect 58578 2 59550 536
rect 59774 2 60746 536
rect 60970 2 61942 536
rect 62166 2 63138 536
rect 63362 2 64242 536
rect 64466 2 65438 536
rect 65662 2 66634 536
rect 66858 2 67830 536
rect 68054 2 69026 536
rect 69250 2 70222 536
rect 70446 2 71418 536
rect 71642 2 72522 536
rect 72746 2 73718 536
rect 73942 2 74914 536
rect 75138 2 76110 536
rect 76334 2 77306 536
rect 77530 2 78502 536
rect 78726 2 79606 536
rect 79830 2 80802 536
rect 81026 2 81998 536
rect 82222 2 83194 536
rect 83418 2 84390 536
rect 84614 2 85586 536
rect 85810 2 86782 536
rect 87006 2 87886 536
rect 88110 2 89082 536
rect 89306 2 90278 536
rect 90502 2 91474 536
rect 91698 2 92670 536
rect 92894 2 93866 536
rect 94090 2 95062 536
rect 95286 2 96166 536
rect 96390 2 97362 536
rect 97586 2 98558 536
rect 98782 2 99754 536
rect 99978 2 100950 536
rect 101174 2 102146 536
rect 102370 2 103250 536
rect 103474 2 104446 536
rect 104670 2 105642 536
rect 105866 2 106838 536
rect 107062 2 108034 536
rect 108258 2 109230 536
rect 109454 2 110426 536
rect 110650 2 111530 536
rect 111754 2 112726 536
rect 112950 2 113922 536
rect 114146 2 115118 536
rect 115342 2 116314 536
rect 116538 2 117510 536
rect 117734 2 118706 536
rect 118930 2 119810 536
rect 120034 2 121006 536
rect 121230 2 122202 536
rect 122426 2 123398 536
rect 123622 2 124594 536
rect 124818 2 125790 536
rect 126014 2 126894 536
rect 127118 2 128090 536
rect 128314 2 129286 536
rect 129510 2 130482 536
rect 130706 2 131678 536
rect 131902 2 132874 536
rect 133098 2 134070 536
rect 134294 2 135174 536
rect 135398 2 136370 536
rect 136594 2 137566 536
rect 137790 2 138762 536
rect 138986 2 139958 536
rect 140182 2 141154 536
rect 141378 2 142350 536
rect 142574 2 143454 536
rect 143678 2 144650 536
rect 144874 2 145846 536
rect 146070 2 147042 536
rect 147266 2 148238 536
rect 148462 2 149434 536
rect 149658 2 150538 536
rect 150762 2 151734 536
rect 151958 2 152930 536
rect 153154 2 154126 536
rect 154350 2 155322 536
rect 155546 2 156518 536
rect 156742 2 157714 536
rect 157938 2 158818 536
rect 159042 2 160014 536
rect 160238 2 161210 536
rect 161434 2 162406 536
rect 162630 2 163602 536
rect 163826 2 164798 536
rect 165022 2 165994 536
rect 166218 2 167098 536
rect 167322 2 168294 536
rect 168518 2 169490 536
rect 169714 2 170686 536
rect 170910 2 171882 536
rect 172106 2 173078 536
rect 173302 2 174182 536
rect 174406 2 175378 536
rect 175602 2 176574 536
rect 176798 2 177770 536
rect 177994 2 178966 536
rect 179190 2 180162 536
rect 180386 2 181358 536
rect 181582 2 182462 536
rect 182686 2 183658 536
rect 183882 2 184854 536
rect 185078 2 186050 536
rect 186274 2 187246 536
rect 187470 2 188442 536
rect 188666 2 189638 536
rect 189862 2 190742 536
rect 190966 2 191938 536
rect 192162 2 193134 536
rect 193358 2 194330 536
rect 194554 2 195526 536
rect 195750 2 196722 536
rect 196946 2 197826 536
rect 198050 2 199022 536
rect 199246 2 200218 536
rect 200442 2 201414 536
rect 201638 2 202610 536
rect 202834 2 203806 536
rect 204030 2 205002 536
rect 205226 2 206106 536
rect 206330 2 207302 536
rect 207526 2 208498 536
rect 208722 2 209694 536
rect 209918 2 210890 536
rect 211114 2 212086 536
rect 212310 2 213282 536
rect 213506 2 214386 536
rect 214610 2 215582 536
rect 215806 2 216778 536
rect 217002 2 217974 536
rect 218198 2 219170 536
rect 219394 2 220366 536
rect 220590 2 221470 536
rect 221694 2 222666 536
rect 222890 2 223862 536
rect 224086 2 225058 536
rect 225282 2 226254 536
rect 226478 2 227450 536
rect 227674 2 228646 536
rect 228870 2 229750 536
rect 229974 2 230946 536
rect 231170 2 232142 536
rect 232366 2 233338 536
rect 233562 2 234534 536
rect 234758 2 235730 536
rect 235954 2 236926 536
rect 237150 2 238030 536
rect 238254 2 239226 536
rect 239450 2 240422 536
rect 240646 2 241618 536
rect 241842 2 242814 536
rect 243038 2 244010 536
rect 244234 2 245114 536
rect 245338 2 246310 536
rect 246534 2 247506 536
rect 247730 2 248702 536
rect 248926 2 249898 536
rect 250122 2 251094 536
rect 251318 2 252290 536
rect 252514 2 253394 536
rect 253618 2 254590 536
rect 254814 2 255786 536
rect 256010 2 256982 536
rect 257206 2 258178 536
rect 258402 2 259374 536
rect 259598 2 260570 536
rect 260794 2 261674 536
rect 261898 2 262870 536
rect 263094 2 264066 536
rect 264290 2 265262 536
rect 265486 2 266458 536
rect 266682 2 267654 536
rect 267878 2 268758 536
rect 268982 2 269954 536
rect 270178 2 271150 536
rect 271374 2 272346 536
rect 272570 2 273542 536
rect 273766 2 274738 536
rect 274962 2 275934 536
rect 276158 2 277038 536
rect 277262 2 278234 536
rect 278458 2 279430 536
rect 279654 2 280626 536
rect 280850 2 281822 536
rect 282046 2 283018 536
rect 283242 2 284214 536
rect 284438 2 285318 536
rect 285542 2 286514 536
rect 286738 2 287710 536
rect 287934 2 288906 536
rect 289130 2 290102 536
rect 290326 2 291298 536
rect 291522 2 292494 536
rect 292718 2 293598 536
rect 293822 2 294794 536
rect 295018 2 295990 536
rect 296214 2 297186 536
rect 297410 2 298382 536
rect 298606 2 299578 536
rect 299802 2 300682 536
rect 300906 2 301878 536
rect 302102 2 303074 536
rect 303298 2 304270 536
rect 304494 2 305466 536
rect 305690 2 306662 536
rect 306886 2 307858 536
rect 308082 2 308962 536
rect 309186 2 310158 536
rect 310382 2 311354 536
rect 311578 2 312550 536
rect 312774 2 313746 536
rect 313970 2 314942 536
rect 315166 2 316138 536
rect 316362 2 317242 536
rect 317466 2 318438 536
rect 318662 2 319634 536
rect 319858 2 320830 536
rect 321054 2 322026 536
rect 322250 2 323222 536
rect 323446 2 324326 536
rect 324550 2 325522 536
rect 325746 2 326718 536
rect 326942 2 327914 536
rect 328138 2 329110 536
rect 329334 2 330306 536
rect 330530 2 331502 536
rect 331726 2 332606 536
rect 332830 2 333802 536
rect 334026 2 334998 536
rect 335222 2 336194 536
rect 336418 2 337390 536
rect 337614 2 338586 536
rect 338810 2 339782 536
rect 340006 2 340886 536
rect 341110 2 342082 536
rect 342306 2 343278 536
rect 343502 2 344474 536
rect 344698 2 345670 536
rect 345894 2 346866 536
rect 347090 2 347970 536
rect 348194 2 349166 536
rect 349390 2 350362 536
rect 350586 2 351558 536
rect 351782 2 352754 536
rect 352978 2 353950 536
rect 354174 2 355146 536
rect 355370 2 356250 536
rect 356474 2 357446 536
rect 357670 2 358642 536
rect 358866 2 359838 536
rect 360062 2 361034 536
rect 361258 2 362230 536
rect 362454 2 363426 536
rect 363650 2 364530 536
rect 364754 2 365726 536
rect 365950 2 366922 536
rect 367146 2 368118 536
rect 368342 2 369314 536
rect 369538 2 370510 536
rect 370734 2 371614 536
rect 371838 2 372810 536
rect 373034 2 374006 536
rect 374230 2 375202 536
rect 375426 2 376398 536
rect 376622 2 377594 536
rect 377818 2 378790 536
rect 379014 2 379894 536
rect 380118 2 381090 536
rect 381314 2 382286 536
rect 382510 2 383482 536
rect 383706 2 384678 536
rect 384902 2 385874 536
rect 386098 2 387070 536
rect 387294 2 388174 536
rect 388398 2 389370 536
rect 389594 2 390566 536
rect 390790 2 391762 536
rect 391986 2 392958 536
rect 393182 2 394154 536
rect 394378 2 395258 536
rect 395482 2 396454 536
rect 396678 2 397650 536
rect 397874 2 398846 536
rect 399070 2 400042 536
rect 400266 2 401238 536
rect 401462 2 402434 536
rect 402658 2 403538 536
rect 403762 2 404734 536
rect 404958 2 405930 536
rect 406154 2 407126 536
rect 407350 2 408322 536
rect 408546 2 409518 536
rect 409742 2 410714 536
rect 410938 2 411818 536
rect 412042 2 413014 536
rect 413238 2 414210 536
rect 414434 2 415406 536
rect 415630 2 416602 536
rect 416826 2 417798 536
rect 418022 2 418902 536
rect 419126 2 420098 536
rect 420322 2 421294 536
rect 421518 2 422490 536
rect 422714 2 423686 536
rect 423910 2 424882 536
rect 425106 2 426078 536
rect 426302 2 427182 536
rect 427406 2 428378 536
rect 428602 2 429574 536
rect 429798 2 430770 536
rect 430994 2 431966 536
rect 432190 2 433162 536
rect 433386 2 434358 536
rect 434582 2 435462 536
rect 435686 2 436658 536
rect 436882 2 437854 536
rect 438078 2 439050 536
rect 439274 2 440246 536
rect 440470 2 441442 536
rect 441666 2 442546 536
rect 442770 2 443742 536
rect 443966 2 444938 536
rect 445162 2 446134 536
rect 446358 2 447330 536
rect 447554 2 448526 536
rect 448750 2 449722 536
rect 449946 2 450826 536
rect 451050 2 452022 536
rect 452246 2 453218 536
rect 453442 2 454414 536
rect 454638 2 455610 536
rect 455834 2 456806 536
rect 457030 2 458002 536
rect 458226 2 459106 536
rect 459330 2 460302 536
rect 460526 2 461498 536
rect 461722 2 462694 536
rect 462918 2 463890 536
rect 464114 2 465086 536
rect 465310 2 466190 536
rect 466414 2 467386 536
rect 467610 2 468582 536
rect 468806 2 469778 536
rect 470002 2 470974 536
rect 471198 2 472170 536
rect 472394 2 473366 536
rect 473590 2 474470 536
rect 474694 2 475666 536
rect 475890 2 476862 536
rect 477086 2 478058 536
rect 478282 2 479254 536
rect 479478 2 480450 536
rect 480674 2 481646 536
rect 481870 2 482750 536
rect 482974 2 483946 536
rect 484170 2 485142 536
rect 485366 2 486338 536
rect 486562 2 487534 536
rect 487758 2 488730 536
rect 488954 2 489834 536
rect 490058 2 491030 536
rect 491254 2 492226 536
rect 492450 2 493422 536
rect 493646 2 494618 536
rect 494842 2 495814 536
rect 496038 2 497010 536
rect 497234 2 498114 536
rect 498338 2 499310 536
rect 499534 2 500506 536
rect 500730 2 501702 536
rect 501926 2 502898 536
rect 503122 2 504094 536
rect 504318 2 505290 536
rect 505514 2 506394 536
rect 506618 2 507590 536
rect 507814 2 508786 536
rect 509010 2 509982 536
rect 510206 2 511178 536
rect 511402 2 512374 536
rect 512598 2 513478 536
rect 513702 2 514674 536
rect 514898 2 515870 536
rect 516094 2 517066 536
rect 517290 2 518262 536
rect 518486 2 519458 536
rect 519682 2 520654 536
rect 520878 2 521758 536
rect 521982 2 522954 536
rect 523178 2 524150 536
rect 524374 2 525346 536
rect 525570 2 526542 536
rect 526766 2 527738 536
rect 527962 2 528934 536
rect 529158 2 530038 536
rect 530262 2 531234 536
rect 531458 2 532430 536
rect 532654 2 533626 536
rect 533850 2 534822 536
rect 535046 2 536018 536
rect 536242 2 537122 536
rect 537346 2 538318 536
rect 538542 2 539514 536
rect 539738 2 540710 536
rect 540934 2 541906 536
rect 542130 2 543102 536
rect 543326 2 544298 536
rect 544522 2 545402 536
rect 545626 2 546598 536
rect 546822 2 547794 536
rect 548018 2 548990 536
rect 549214 2 550186 536
rect 550410 2 551382 536
rect 551606 2 552578 536
rect 552802 2 553682 536
rect 553906 2 554878 536
rect 555102 2 556074 536
rect 556298 2 557270 536
rect 557494 2 558466 536
rect 558690 2 559662 536
rect 559886 2 560766 536
rect 560990 2 561962 536
rect 562186 2 563158 536
rect 563382 2 564354 536
rect 564578 2 565550 536
rect 565774 2 566746 536
rect 566970 2 567942 536
rect 568166 2 569046 536
rect 569270 2 570242 536
rect 570466 2 571438 536
rect 571662 2 572634 536
rect 572858 2 573830 536
rect 574054 2 575026 536
rect 575250 2 576222 536
rect 576446 2 577326 536
rect 577550 2 578522 536
rect 578746 2 579718 536
rect 579942 2 580914 536
rect 581138 2 582110 536
rect 582334 2 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 105 189036 578943 189141
rect 560 188636 578943 189036
rect 105 176116 578943 188636
rect 560 175716 578943 176116
rect 105 163060 578943 175716
rect 560 162660 578943 163060
rect 105 150004 578943 162660
rect 560 149604 578943 150004
rect 105 136948 578943 149604
rect 560 136548 578943 136948
rect 105 123892 578943 136548
rect 560 123492 578943 123892
rect 105 110836 578943 123492
rect 560 110436 578943 110836
rect 105 97780 578943 110436
rect 560 97380 578943 97780
rect 105 84860 578943 97380
rect 560 84460 578943 84860
rect 105 71804 578943 84460
rect 560 71404 578943 71804
rect 105 58748 578943 71404
rect 560 58348 578943 58748
rect 105 45692 578943 58348
rect 560 45292 578943 45692
rect 105 32636 578943 45292
rect 560 32236 578943 32636
rect 105 19580 578943 32236
rect 560 19180 578943 19580
rect 105 6660 578943 19180
rect 560 6260 578943 6660
rect 105 443 578943 6260
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -1894 2414 705830
rect 5514 -3814 6134 707750
rect 9234 106800 9854 709670
rect 12954 193500 13574 711590
rect 19794 193500 20414 705830
rect 23514 193500 24134 707750
rect 27234 193500 27854 709670
rect 30954 193500 31574 711590
rect 37794 193500 38414 705830
rect 41514 193500 42134 707750
rect 45234 193500 45854 709670
rect 48954 193500 49574 711590
rect 55794 193500 56414 705830
rect 59514 193500 60134 707750
rect 63234 193500 63854 709670
rect 66954 193500 67574 711590
rect 73794 193500 74414 705830
rect 77514 193500 78134 707750
rect 81234 193500 81854 709670
rect 84954 193500 85574 711590
rect 91794 193500 92414 705830
rect 95514 193500 96134 707750
rect 99234 193500 99854 709670
rect 102954 193500 103574 711590
rect 109794 193500 110414 705830
rect 113514 193500 114134 707750
rect 117234 193500 117854 709670
rect 120954 193500 121574 711590
rect 127794 107308 128414 705830
rect 131514 107308 132134 707750
rect 135234 107308 135854 709670
rect 138954 107308 139574 711590
rect 145794 107308 146414 705830
rect 149514 107308 150134 707750
rect 153234 107308 153854 709670
rect 156954 107308 157574 711590
rect 163794 107308 164414 705830
rect 167514 107308 168134 707750
rect 171234 107308 171854 709670
rect 174954 107308 175574 711590
rect 181794 107308 182414 705830
rect 185514 107308 186134 707750
rect 189234 107308 189854 709670
rect 192954 107308 193574 711590
rect 199794 107308 200414 705830
rect 203514 107308 204134 707750
rect 207234 107308 207854 709670
rect 210954 107308 211574 711590
rect 217794 107308 218414 705830
rect 221514 107308 222134 707750
rect 225234 107308 225854 709670
rect 228954 107308 229574 711590
rect 235794 107308 236414 705830
rect 239514 107308 240134 707750
rect 243234 107308 243854 709670
rect 246954 107308 247574 711590
rect 9234 -5734 9854 4000
rect 12954 -7654 13574 4000
rect 19794 -1894 20414 4000
rect 23514 -3814 24134 4000
rect 27234 -5734 27854 4000
rect 30954 -7654 31574 4000
rect 37794 -1894 38414 4000
rect 41514 -3814 42134 4000
rect 45234 -5734 45854 4000
rect 48954 -7654 49574 4000
rect 55794 -1894 56414 4000
rect 59514 -3814 60134 4000
rect 63234 -5734 63854 4000
rect 66954 -7654 67574 4000
rect 73794 -1894 74414 4000
rect 77514 -3814 78134 4000
rect 81234 -5734 81854 4000
rect 84954 -7654 85574 4000
rect 91794 -1894 92414 4000
rect 95514 -3814 96134 4000
rect 99234 -5734 99854 4000
rect 102954 -7654 103574 4000
rect 109794 -1894 110414 4000
rect 113514 -3814 114134 4000
rect 117234 -5734 117854 4000
rect 120954 -7654 121574 4000
rect 127794 -1894 128414 4000
rect 131514 -3814 132134 4000
rect 135234 -5734 135854 4000
rect 138954 -7654 139574 4000
rect 145794 -1894 146414 4000
rect 149514 -3814 150134 4000
rect 153234 -5734 153854 4000
rect 156954 -7654 157574 4000
rect 163794 -1894 164414 4000
rect 167514 -3814 168134 4000
rect 171234 -5734 171854 4000
rect 174954 -7654 175574 4000
rect 181794 -1894 182414 4000
rect 185514 -3814 186134 4000
rect 189234 -5734 189854 4000
rect 192954 -7654 193574 4000
rect 199794 -1894 200414 4000
rect 203514 -3814 204134 4000
rect 207234 -5734 207854 4000
rect 210954 -7654 211574 4000
rect 217794 -1894 218414 4000
rect 221514 -3814 222134 4000
rect 225234 -5734 225854 4000
rect 228954 -7654 229574 4000
rect 235794 -1894 236414 4000
rect 239514 -3814 240134 4000
rect 243234 -5734 243854 4000
rect 246954 -7654 247574 4000
rect 253794 -1894 254414 705830
rect 257514 -3814 258134 707750
rect 261234 -5734 261854 709670
rect 264954 -7654 265574 711590
rect 271794 -1894 272414 705830
rect 275514 -3814 276134 707750
rect 279234 -5734 279854 709670
rect 282954 -7654 283574 711590
rect 289794 -1894 290414 705830
rect 293514 -3814 294134 707750
rect 297234 -5734 297854 709670
rect 300954 -7654 301574 711590
rect 307794 -1894 308414 705830
rect 311514 -3814 312134 707750
rect 315234 -5734 315854 709670
rect 318954 -7654 319574 711590
rect 325794 -1894 326414 705830
rect 329514 -3814 330134 707750
rect 333234 -5734 333854 709670
rect 336954 -7654 337574 711590
rect 343794 -1894 344414 705830
rect 347514 -3814 348134 707750
rect 351234 -5734 351854 709670
rect 354954 -7654 355574 711590
rect 361794 -1894 362414 705830
rect 365514 -3814 366134 707750
rect 369234 -5734 369854 709670
rect 372954 -7654 373574 711590
rect 379794 -1894 380414 705830
rect 383514 -3814 384134 707750
rect 387234 -5734 387854 709670
rect 390954 -7654 391574 711590
rect 397794 -1894 398414 705830
rect 401514 -3814 402134 707750
rect 405234 -5734 405854 709670
rect 408954 -7654 409574 711590
rect 415794 -1894 416414 705830
rect 419514 -3814 420134 707750
rect 423234 -5734 423854 709670
rect 426954 -7654 427574 711590
rect 433794 -1894 434414 705830
rect 437514 -3814 438134 707750
rect 441234 -5734 441854 709670
rect 444954 -7654 445574 711590
rect 451794 -1894 452414 705830
rect 455514 -3814 456134 707750
rect 459234 -5734 459854 709670
rect 462954 -7654 463574 711590
rect 469794 -1894 470414 705830
rect 473514 -3814 474134 707750
rect 477234 -5734 477854 709670
rect 480954 -7654 481574 711590
rect 487794 -1894 488414 705830
rect 491514 -3814 492134 707750
rect 495234 -5734 495854 709670
rect 498954 -7654 499574 711590
rect 505794 -1894 506414 705830
rect 509514 -3814 510134 707750
rect 513234 -5734 513854 709670
rect 516954 -7654 517574 711590
rect 523794 -1894 524414 705830
rect 527514 -3814 528134 707750
rect 531234 -5734 531854 709670
rect 534954 -7654 535574 711590
rect 541794 -1894 542414 705830
rect 545514 -3814 546134 707750
rect 549234 -5734 549854 709670
rect 552954 -7654 553574 711590
rect 559794 -1894 560414 705830
rect 563514 -3814 564134 707750
rect 567234 -5734 567854 709670
rect 570954 -7654 571574 711590
rect 577794 -1894 578414 705830
rect 581514 -3814 582134 707750
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 12203 107228 127714 188053
rect 128494 107228 131434 188053
rect 132214 107228 135154 188053
rect 135934 107228 138874 188053
rect 139654 107228 145714 188053
rect 146494 107228 149434 188053
rect 150214 107228 153154 188053
rect 153934 107228 156874 188053
rect 157654 107228 163714 188053
rect 164494 107228 167434 188053
rect 168214 107228 171154 188053
rect 171934 107228 174874 188053
rect 175654 107228 181714 188053
rect 182494 107228 185434 188053
rect 186214 107228 189154 188053
rect 189934 107228 192874 188053
rect 193654 107228 199714 188053
rect 200494 107228 203434 188053
rect 204214 107228 207154 188053
rect 207934 107228 210874 188053
rect 211654 107228 217714 188053
rect 218494 107228 221434 188053
rect 222214 107228 225154 188053
rect 225934 107228 228874 188053
rect 229654 107228 235714 188053
rect 236494 107228 239434 188053
rect 240214 107228 240245 188053
rect 12203 4080 240245 107228
rect 12203 715 12874 4080
rect 13654 715 19714 4080
rect 20494 715 23434 4080
rect 24214 715 27154 4080
rect 27934 715 30874 4080
rect 31654 715 37714 4080
rect 38494 715 41434 4080
rect 42214 715 45154 4080
rect 45934 715 48874 4080
rect 49654 715 55714 4080
rect 56494 715 59434 4080
rect 60214 715 63154 4080
rect 63934 715 66874 4080
rect 67654 715 73714 4080
rect 74494 715 77434 4080
rect 78214 715 81154 4080
rect 81934 715 84874 4080
rect 85654 715 91714 4080
rect 92494 715 95434 4080
rect 96214 715 99154 4080
rect 99934 715 102874 4080
rect 103654 715 109714 4080
rect 110494 715 113434 4080
rect 114214 715 117154 4080
rect 117934 715 120874 4080
rect 121654 715 127714 4080
rect 128494 715 131434 4080
rect 132214 715 135154 4080
rect 135934 715 138874 4080
rect 139654 715 145714 4080
rect 146494 715 149434 4080
rect 150214 715 153154 4080
rect 153934 715 156874 4080
rect 157654 715 163714 4080
rect 164494 715 167434 4080
rect 168214 715 171154 4080
rect 171934 715 174874 4080
rect 175654 715 181714 4080
rect 182494 715 185434 4080
rect 186214 715 189154 4080
rect 189934 715 192874 4080
rect 193654 715 199714 4080
rect 200494 715 203434 4080
rect 204214 715 207154 4080
rect 207934 715 210874 4080
rect 211654 715 217714 4080
rect 218494 715 221434 4080
rect 222214 715 225154 4080
rect 225934 715 228874 4080
rect 229654 715 235714 4080
rect 236494 715 239434 4080
rect 240214 715 240245 4080
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 698026 592650 698646
rect -6806 694306 590730 694926
rect -4886 690586 588810 691206
rect -2966 686866 586890 687486
rect -8726 680026 592650 680646
rect -6806 676306 590730 676926
rect -4886 672586 588810 673206
rect -2966 668866 586890 669486
rect -8726 662026 592650 662646
rect -6806 658306 590730 658926
rect -4886 654586 588810 655206
rect -2966 650866 586890 651486
rect -8726 644026 592650 644646
rect -6806 640306 590730 640926
rect -4886 636586 588810 637206
rect -2966 632866 586890 633486
rect -8726 626026 592650 626646
rect -6806 622306 590730 622926
rect -4886 618586 588810 619206
rect -2966 614866 586890 615486
rect -8726 608026 592650 608646
rect -6806 604306 590730 604926
rect -4886 600586 588810 601206
rect -2966 596866 586890 597486
rect -8726 590026 592650 590646
rect -6806 586306 590730 586926
rect -4886 582586 588810 583206
rect -2966 578866 586890 579486
rect -8726 572026 592650 572646
rect -6806 568306 590730 568926
rect -4886 564586 588810 565206
rect -2966 560866 586890 561486
rect -8726 554026 592650 554646
rect -6806 550306 590730 550926
rect -4886 546586 588810 547206
rect -2966 542866 586890 543486
rect -8726 536026 592650 536646
rect -6806 532306 590730 532926
rect -4886 528586 588810 529206
rect -2966 524866 586890 525486
rect -8726 518026 592650 518646
rect -6806 514306 590730 514926
rect -4886 510586 588810 511206
rect -2966 506866 586890 507486
rect -8726 500026 592650 500646
rect -6806 496306 590730 496926
rect -4886 492586 588810 493206
rect -2966 488866 586890 489486
rect -8726 482026 592650 482646
rect -6806 478306 590730 478926
rect -4886 474586 588810 475206
rect -2966 470866 586890 471486
rect -8726 464026 592650 464646
rect -6806 460306 590730 460926
rect -4886 456586 588810 457206
rect -2966 452866 586890 453486
rect -8726 446026 592650 446646
rect -6806 442306 590730 442926
rect -4886 438586 588810 439206
rect -2966 434866 586890 435486
rect -8726 428026 592650 428646
rect -6806 424306 590730 424926
rect -4886 420586 588810 421206
rect -2966 416866 586890 417486
rect -8726 410026 592650 410646
rect -6806 406306 590730 406926
rect -4886 402586 588810 403206
rect -2966 398866 586890 399486
rect -8726 392026 592650 392646
rect -6806 388306 590730 388926
rect -4886 384586 588810 385206
rect -2966 380866 586890 381486
rect -8726 374026 592650 374646
rect -6806 370306 590730 370926
rect -4886 366586 588810 367206
rect -2966 362866 586890 363486
rect -8726 356026 592650 356646
rect -6806 352306 590730 352926
rect -4886 348586 588810 349206
rect -2966 344866 586890 345486
rect -8726 338026 592650 338646
rect -6806 334306 590730 334926
rect -4886 330586 588810 331206
rect -2966 326866 586890 327486
rect -8726 320026 592650 320646
rect -6806 316306 590730 316926
rect -4886 312586 588810 313206
rect -2966 308866 586890 309486
rect -8726 302026 592650 302646
rect -6806 298306 590730 298926
rect -4886 294586 588810 295206
rect -2966 290866 586890 291486
rect -8726 284026 592650 284646
rect -6806 280306 590730 280926
rect -4886 276586 588810 277206
rect -2966 272866 586890 273486
rect -8726 266026 592650 266646
rect -6806 262306 590730 262926
rect -4886 258586 588810 259206
rect -2966 254866 586890 255486
rect -8726 248026 592650 248646
rect -6806 244306 590730 244926
rect -4886 240586 588810 241206
rect -2966 236866 586890 237486
rect -8726 230026 592650 230646
rect -6806 226306 590730 226926
rect -4886 222586 588810 223206
rect -2966 218866 586890 219486
rect -8726 212026 592650 212646
rect -6806 208306 590730 208926
rect -4886 204586 588810 205206
rect -2966 200866 586890 201486
rect -8726 194026 592650 194646
rect -6806 190306 590730 190926
rect -4886 186586 588810 187206
rect -2966 182866 586890 183486
rect -8726 176026 592650 176646
rect -6806 172306 590730 172926
rect -4886 168586 588810 169206
rect -2966 164866 586890 165486
rect -8726 158026 592650 158646
rect -6806 154306 590730 154926
rect -4886 150586 588810 151206
rect -2966 146866 586890 147486
rect -8726 140026 592650 140646
rect -6806 136306 590730 136926
rect -4886 132586 588810 133206
rect -2966 128866 586890 129486
rect -8726 122026 592650 122646
rect -6806 118306 590730 118926
rect -4886 114586 588810 115206
rect -2966 110866 586890 111486
rect -8726 104026 592650 104646
rect -6806 100306 590730 100926
rect -4886 96586 588810 97206
rect -2966 92866 586890 93486
rect -8726 86026 592650 86646
rect -6806 82306 590730 82926
rect -4886 78586 588810 79206
rect -2966 74866 586890 75486
rect -8726 68026 592650 68646
rect -6806 64306 590730 64926
rect -4886 60586 588810 61206
rect -2966 56866 586890 57486
rect -8726 50026 592650 50646
rect -6806 46306 590730 46926
rect -4886 42586 588810 43206
rect -2966 38866 586890 39486
rect -8726 32026 592650 32646
rect -6806 28306 590730 28926
rect -4886 24586 588810 25206
rect -2966 20866 586890 21486
rect -8726 14026 592650 14646
rect -6806 10306 590730 10926
rect -4886 6586 588810 7206
rect -2966 2866 586890 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 532 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 -1894 38414 4000 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 -1894 74414 4000 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 -1894 110414 4000 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 -1894 146414 4000 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 -1894 182414 4000 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 -1894 218414 4000 6 vccd1
port 532 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 37794 193500 38414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 73794 193500 74414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 109794 193500 110414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 145794 107308 146414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 181794 107308 182414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 217794 107308 218414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 532 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 532 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 533 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 533 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 41514 -3814 42134 4000 6 vccd2
port 533 nsew power input
rlabel metal4 s 77514 -3814 78134 4000 6 vccd2
port 533 nsew power input
rlabel metal4 s 113514 -3814 114134 4000 6 vccd2
port 533 nsew power input
rlabel metal4 s 149514 -3814 150134 4000 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 -3814 186134 4000 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 -3814 222134 4000 6 vccd2
port 533 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 41514 193500 42134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 77514 193500 78134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 113514 193500 114134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 149514 107308 150134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 185514 107308 186134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 221514 107308 222134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 533 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 533 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 534 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 534 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 9234 -5734 9854 4000 8 vdda1
port 534 nsew power input
rlabel metal4 s 45234 -5734 45854 4000 8 vdda1
port 534 nsew power input
rlabel metal4 s 81234 -5734 81854 4000 8 vdda1
port 534 nsew power input
rlabel metal4 s 117234 -5734 117854 4000 8 vdda1
port 534 nsew power input
rlabel metal4 s 153234 -5734 153854 4000 8 vdda1
port 534 nsew power input
rlabel metal4 s 189234 -5734 189854 4000 8 vdda1
port 534 nsew power input
rlabel metal4 s 225234 -5734 225854 4000 8 vdda1
port 534 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power input
rlabel metal4 s 9234 106800 9854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 45234 193500 45854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 81234 193500 81854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 117234 193500 117854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 153234 107308 153854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 189234 107308 189854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 225234 107308 225854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 534 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 534 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 535 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 535 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 12954 -7654 13574 4000 8 vdda2
port 535 nsew power input
rlabel metal4 s 48954 -7654 49574 4000 8 vdda2
port 535 nsew power input
rlabel metal4 s 84954 -7654 85574 4000 8 vdda2
port 535 nsew power input
rlabel metal4 s 120954 -7654 121574 4000 8 vdda2
port 535 nsew power input
rlabel metal4 s 156954 -7654 157574 4000 8 vdda2
port 535 nsew power input
rlabel metal4 s 192954 -7654 193574 4000 8 vdda2
port 535 nsew power input
rlabel metal4 s 228954 -7654 229574 4000 8 vdda2
port 535 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power input
rlabel metal4 s 12954 193500 13574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 48954 193500 49574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 84954 193500 85574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 120954 193500 121574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 156954 107308 157574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 192954 107308 193574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 228954 107308 229574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 535 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 535 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 536 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 27234 -5734 27854 4000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 63234 -5734 63854 4000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 -5734 99854 4000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 -5734 135854 4000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 171234 -5734 171854 4000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 207234 -5734 207854 4000 8 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 -5734 243854 4000 8 vssa1
port 536 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground input
rlabel metal4 s 27234 193500 27854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 63234 193500 63854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 99234 193500 99854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 135234 107308 135854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 171234 107308 171854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 207234 107308 207854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 243234 107308 243854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 536 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 537 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 30954 -7654 31574 4000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 66954 -7654 67574 4000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 -7654 103574 4000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 -7654 139574 4000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 174954 -7654 175574 4000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 210954 -7654 211574 4000 8 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 -7654 247574 4000 8 vssa2
port 537 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground input
rlabel metal4 s 30954 193500 31574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 66954 193500 67574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 102954 193500 103574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 138954 107308 139574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 174954 107308 175574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 210954 107308 211574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 246954 107308 247574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 537 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 538 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 19794 -1894 20414 4000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 55794 -1894 56414 4000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 -1894 92414 4000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 -1894 128414 4000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 163794 -1894 164414 4000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 199794 -1894 200414 4000 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 -1894 236414 4000 6 vssd1
port 538 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground input
rlabel metal4 s 19794 193500 20414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 55794 193500 56414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 91794 193500 92414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 127794 107308 128414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 163794 107308 164414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 199794 107308 200414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 235794 107308 236414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 538 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 539 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 23514 -3814 24134 4000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 59514 -3814 60134 4000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 -3814 96134 4000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 -3814 132134 4000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 167514 -3814 168134 4000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 203514 -3814 204134 4000 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 -3814 240134 4000 6 vssd2
port 539 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground input
rlabel metal4 s 23514 193500 24134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 59514 193500 60134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 95514 193500 96134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 131514 107308 132134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 167514 107308 168134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 203514 107308 204134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 239514 107308 240134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 539 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 48165892
string GDS_FILE /home/re19/Caravel/temporal_runtime_monitor/openlane/user_project_wrapper/runs/user_project_wrapper/results/finishing/user_project_wrapper.magic.gds
string GDS_START 46582784
<< end >>

