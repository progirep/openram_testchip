magic
tech sky130A
magscale 1 2
timestamp 1646995934
<< obsli1 >>
rect 1104 2159 238832 117521
<< obsm1 >>
rect 750 1844 239186 117552
<< metal2 >>
rect 754 119200 810 120000
rect 2318 119200 2374 120000
rect 3974 119200 4030 120000
rect 5538 119200 5594 120000
rect 7194 119200 7250 120000
rect 8758 119200 8814 120000
rect 10414 119200 10470 120000
rect 11978 119200 12034 120000
rect 13634 119200 13690 120000
rect 15198 119200 15254 120000
rect 16854 119200 16910 120000
rect 18418 119200 18474 120000
rect 20074 119200 20130 120000
rect 21638 119200 21694 120000
rect 23294 119200 23350 120000
rect 24858 119200 24914 120000
rect 26514 119200 26570 120000
rect 28078 119200 28134 120000
rect 29734 119200 29790 120000
rect 31298 119200 31354 120000
rect 32954 119200 33010 120000
rect 34518 119200 34574 120000
rect 36174 119200 36230 120000
rect 37738 119200 37794 120000
rect 39394 119200 39450 120000
rect 40958 119200 41014 120000
rect 42614 119200 42670 120000
rect 44178 119200 44234 120000
rect 45834 119200 45890 120000
rect 47398 119200 47454 120000
rect 49054 119200 49110 120000
rect 50618 119200 50674 120000
rect 52274 119200 52330 120000
rect 53838 119200 53894 120000
rect 55494 119200 55550 120000
rect 57058 119200 57114 120000
rect 58714 119200 58770 120000
rect 60278 119200 60334 120000
rect 61934 119200 61990 120000
rect 63498 119200 63554 120000
rect 65154 119200 65210 120000
rect 66718 119200 66774 120000
rect 68374 119200 68430 120000
rect 69938 119200 69994 120000
rect 71594 119200 71650 120000
rect 73158 119200 73214 120000
rect 74814 119200 74870 120000
rect 76378 119200 76434 120000
rect 78034 119200 78090 120000
rect 79598 119200 79654 120000
rect 81254 119200 81310 120000
rect 82910 119200 82966 120000
rect 84474 119200 84530 120000
rect 86130 119200 86186 120000
rect 87694 119200 87750 120000
rect 89350 119200 89406 120000
rect 90914 119200 90970 120000
rect 92570 119200 92626 120000
rect 94134 119200 94190 120000
rect 95790 119200 95846 120000
rect 97354 119200 97410 120000
rect 99010 119200 99066 120000
rect 100574 119200 100630 120000
rect 102230 119200 102286 120000
rect 103794 119200 103850 120000
rect 105450 119200 105506 120000
rect 107014 119200 107070 120000
rect 108670 119200 108726 120000
rect 110234 119200 110290 120000
rect 111890 119200 111946 120000
rect 113454 119200 113510 120000
rect 115110 119200 115166 120000
rect 116674 119200 116730 120000
rect 118330 119200 118386 120000
rect 119894 119200 119950 120000
rect 121550 119200 121606 120000
rect 123114 119200 123170 120000
rect 124770 119200 124826 120000
rect 126334 119200 126390 120000
rect 127990 119200 128046 120000
rect 129554 119200 129610 120000
rect 131210 119200 131266 120000
rect 132774 119200 132830 120000
rect 134430 119200 134486 120000
rect 135994 119200 136050 120000
rect 137650 119200 137706 120000
rect 139214 119200 139270 120000
rect 140870 119200 140926 120000
rect 142434 119200 142490 120000
rect 144090 119200 144146 120000
rect 145654 119200 145710 120000
rect 147310 119200 147366 120000
rect 148874 119200 148930 120000
rect 150530 119200 150586 120000
rect 152094 119200 152150 120000
rect 153750 119200 153806 120000
rect 155314 119200 155370 120000
rect 156970 119200 157026 120000
rect 158534 119200 158590 120000
rect 160190 119200 160246 120000
rect 161846 119200 161902 120000
rect 163410 119200 163466 120000
rect 165066 119200 165122 120000
rect 166630 119200 166686 120000
rect 168286 119200 168342 120000
rect 169850 119200 169906 120000
rect 171506 119200 171562 120000
rect 173070 119200 173126 120000
rect 174726 119200 174782 120000
rect 176290 119200 176346 120000
rect 177946 119200 178002 120000
rect 179510 119200 179566 120000
rect 181166 119200 181222 120000
rect 182730 119200 182786 120000
rect 184386 119200 184442 120000
rect 185950 119200 186006 120000
rect 187606 119200 187662 120000
rect 189170 119200 189226 120000
rect 190826 119200 190882 120000
rect 192390 119200 192446 120000
rect 194046 119200 194102 120000
rect 195610 119200 195666 120000
rect 197266 119200 197322 120000
rect 198830 119200 198886 120000
rect 200486 119200 200542 120000
rect 202050 119200 202106 120000
rect 203706 119200 203762 120000
rect 205270 119200 205326 120000
rect 206926 119200 206982 120000
rect 208490 119200 208546 120000
rect 210146 119200 210202 120000
rect 211710 119200 211766 120000
rect 213366 119200 213422 120000
rect 214930 119200 214986 120000
rect 216586 119200 216642 120000
rect 218150 119200 218206 120000
rect 219806 119200 219862 120000
rect 221370 119200 221426 120000
rect 223026 119200 223082 120000
rect 224590 119200 224646 120000
rect 226246 119200 226302 120000
rect 227810 119200 227866 120000
rect 229466 119200 229522 120000
rect 231030 119200 231086 120000
rect 232686 119200 232742 120000
rect 234250 119200 234306 120000
rect 235906 119200 235962 120000
rect 237470 119200 237526 120000
rect 239126 119200 239182 120000
rect 846 0 902 800
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5814 0 5870 800
rect 7470 0 7526 800
rect 9218 0 9274 800
rect 10874 0 10930 800
rect 12530 0 12586 800
rect 14186 0 14242 800
rect 15934 0 15990 800
rect 17590 0 17646 800
rect 19246 0 19302 800
rect 20902 0 20958 800
rect 22650 0 22706 800
rect 24306 0 24362 800
rect 25962 0 26018 800
rect 27618 0 27674 800
rect 29366 0 29422 800
rect 31022 0 31078 800
rect 32678 0 32734 800
rect 34334 0 34390 800
rect 36082 0 36138 800
rect 37738 0 37794 800
rect 39394 0 39450 800
rect 41050 0 41106 800
rect 42798 0 42854 800
rect 44454 0 44510 800
rect 46110 0 46166 800
rect 47766 0 47822 800
rect 49514 0 49570 800
rect 51170 0 51226 800
rect 52826 0 52882 800
rect 54482 0 54538 800
rect 56230 0 56286 800
rect 57886 0 57942 800
rect 59542 0 59598 800
rect 61198 0 61254 800
rect 62946 0 63002 800
rect 64602 0 64658 800
rect 66258 0 66314 800
rect 67914 0 67970 800
rect 69662 0 69718 800
rect 71318 0 71374 800
rect 72974 0 73030 800
rect 74630 0 74686 800
rect 76378 0 76434 800
rect 78034 0 78090 800
rect 79690 0 79746 800
rect 81346 0 81402 800
rect 83002 0 83058 800
rect 84750 0 84806 800
rect 86406 0 86462 800
rect 88062 0 88118 800
rect 89718 0 89774 800
rect 91466 0 91522 800
rect 93122 0 93178 800
rect 94778 0 94834 800
rect 96434 0 96490 800
rect 98182 0 98238 800
rect 99838 0 99894 800
rect 101494 0 101550 800
rect 103150 0 103206 800
rect 104898 0 104954 800
rect 106554 0 106610 800
rect 108210 0 108266 800
rect 109866 0 109922 800
rect 111614 0 111670 800
rect 113270 0 113326 800
rect 114926 0 114982 800
rect 116582 0 116638 800
rect 118330 0 118386 800
rect 119986 0 120042 800
rect 121642 0 121698 800
rect 123298 0 123354 800
rect 125046 0 125102 800
rect 126702 0 126758 800
rect 128358 0 128414 800
rect 130014 0 130070 800
rect 131762 0 131818 800
rect 133418 0 133474 800
rect 135074 0 135130 800
rect 136730 0 136786 800
rect 138478 0 138534 800
rect 140134 0 140190 800
rect 141790 0 141846 800
rect 143446 0 143502 800
rect 145194 0 145250 800
rect 146850 0 146906 800
rect 148506 0 148562 800
rect 150162 0 150218 800
rect 151910 0 151966 800
rect 153566 0 153622 800
rect 155222 0 155278 800
rect 156878 0 156934 800
rect 158626 0 158682 800
rect 160282 0 160338 800
rect 161938 0 161994 800
rect 163594 0 163650 800
rect 165250 0 165306 800
rect 166998 0 167054 800
rect 168654 0 168710 800
rect 170310 0 170366 800
rect 171966 0 172022 800
rect 173714 0 173770 800
rect 175370 0 175426 800
rect 177026 0 177082 800
rect 178682 0 178738 800
rect 180430 0 180486 800
rect 182086 0 182142 800
rect 183742 0 183798 800
rect 185398 0 185454 800
rect 187146 0 187202 800
rect 188802 0 188858 800
rect 190458 0 190514 800
rect 192114 0 192170 800
rect 193862 0 193918 800
rect 195518 0 195574 800
rect 197174 0 197230 800
rect 198830 0 198886 800
rect 200578 0 200634 800
rect 202234 0 202290 800
rect 203890 0 203946 800
rect 205546 0 205602 800
rect 207294 0 207350 800
rect 208950 0 209006 800
rect 210606 0 210662 800
rect 212262 0 212318 800
rect 214010 0 214066 800
rect 215666 0 215722 800
rect 217322 0 217378 800
rect 218978 0 219034 800
rect 220726 0 220782 800
rect 222382 0 222438 800
rect 224038 0 224094 800
rect 225694 0 225750 800
rect 227442 0 227498 800
rect 229098 0 229154 800
rect 230754 0 230810 800
rect 232410 0 232466 800
rect 234158 0 234214 800
rect 235814 0 235870 800
rect 237470 0 237526 800
rect 239126 0 239182 800
<< obsm2 >>
rect 866 119144 2262 119354
rect 2430 119144 3918 119354
rect 4086 119144 5482 119354
rect 5650 119144 7138 119354
rect 7306 119144 8702 119354
rect 8870 119144 10358 119354
rect 10526 119144 11922 119354
rect 12090 119144 13578 119354
rect 13746 119144 15142 119354
rect 15310 119144 16798 119354
rect 16966 119144 18362 119354
rect 18530 119144 20018 119354
rect 20186 119144 21582 119354
rect 21750 119144 23238 119354
rect 23406 119144 24802 119354
rect 24970 119144 26458 119354
rect 26626 119144 28022 119354
rect 28190 119144 29678 119354
rect 29846 119144 31242 119354
rect 31410 119144 32898 119354
rect 33066 119144 34462 119354
rect 34630 119144 36118 119354
rect 36286 119144 37682 119354
rect 37850 119144 39338 119354
rect 39506 119144 40902 119354
rect 41070 119144 42558 119354
rect 42726 119144 44122 119354
rect 44290 119144 45778 119354
rect 45946 119144 47342 119354
rect 47510 119144 48998 119354
rect 49166 119144 50562 119354
rect 50730 119144 52218 119354
rect 52386 119144 53782 119354
rect 53950 119144 55438 119354
rect 55606 119144 57002 119354
rect 57170 119144 58658 119354
rect 58826 119144 60222 119354
rect 60390 119144 61878 119354
rect 62046 119144 63442 119354
rect 63610 119144 65098 119354
rect 65266 119144 66662 119354
rect 66830 119144 68318 119354
rect 68486 119144 69882 119354
rect 70050 119144 71538 119354
rect 71706 119144 73102 119354
rect 73270 119144 74758 119354
rect 74926 119144 76322 119354
rect 76490 119144 77978 119354
rect 78146 119144 79542 119354
rect 79710 119144 81198 119354
rect 81366 119144 82854 119354
rect 83022 119144 84418 119354
rect 84586 119144 86074 119354
rect 86242 119144 87638 119354
rect 87806 119144 89294 119354
rect 89462 119144 90858 119354
rect 91026 119144 92514 119354
rect 92682 119144 94078 119354
rect 94246 119144 95734 119354
rect 95902 119144 97298 119354
rect 97466 119144 98954 119354
rect 99122 119144 100518 119354
rect 100686 119144 102174 119354
rect 102342 119144 103738 119354
rect 103906 119144 105394 119354
rect 105562 119144 106958 119354
rect 107126 119144 108614 119354
rect 108782 119144 110178 119354
rect 110346 119144 111834 119354
rect 112002 119144 113398 119354
rect 113566 119144 115054 119354
rect 115222 119144 116618 119354
rect 116786 119144 118274 119354
rect 118442 119144 119838 119354
rect 120006 119144 121494 119354
rect 121662 119144 123058 119354
rect 123226 119144 124714 119354
rect 124882 119144 126278 119354
rect 126446 119144 127934 119354
rect 128102 119144 129498 119354
rect 129666 119144 131154 119354
rect 131322 119144 132718 119354
rect 132886 119144 134374 119354
rect 134542 119144 135938 119354
rect 136106 119144 137594 119354
rect 137762 119144 139158 119354
rect 139326 119144 140814 119354
rect 140982 119144 142378 119354
rect 142546 119144 144034 119354
rect 144202 119144 145598 119354
rect 145766 119144 147254 119354
rect 147422 119144 148818 119354
rect 148986 119144 150474 119354
rect 150642 119144 152038 119354
rect 152206 119144 153694 119354
rect 153862 119144 155258 119354
rect 155426 119144 156914 119354
rect 157082 119144 158478 119354
rect 158646 119144 160134 119354
rect 160302 119144 161790 119354
rect 161958 119144 163354 119354
rect 163522 119144 165010 119354
rect 165178 119144 166574 119354
rect 166742 119144 168230 119354
rect 168398 119144 169794 119354
rect 169962 119144 171450 119354
rect 171618 119144 173014 119354
rect 173182 119144 174670 119354
rect 174838 119144 176234 119354
rect 176402 119144 177890 119354
rect 178058 119144 179454 119354
rect 179622 119144 181110 119354
rect 181278 119144 182674 119354
rect 182842 119144 184330 119354
rect 184498 119144 185894 119354
rect 186062 119144 187550 119354
rect 187718 119144 189114 119354
rect 189282 119144 190770 119354
rect 190938 119144 192334 119354
rect 192502 119144 193990 119354
rect 194158 119144 195554 119354
rect 195722 119144 197210 119354
rect 197378 119144 198774 119354
rect 198942 119144 200430 119354
rect 200598 119144 201994 119354
rect 202162 119144 203650 119354
rect 203818 119144 205214 119354
rect 205382 119144 206870 119354
rect 207038 119144 208434 119354
rect 208602 119144 210090 119354
rect 210258 119144 211654 119354
rect 211822 119144 213310 119354
rect 213478 119144 214874 119354
rect 215042 119144 216530 119354
rect 216698 119144 218094 119354
rect 218262 119144 219750 119354
rect 219918 119144 221314 119354
rect 221482 119144 222970 119354
rect 223138 119144 224534 119354
rect 224702 119144 226190 119354
rect 226358 119144 227754 119354
rect 227922 119144 229410 119354
rect 229578 119144 230974 119354
rect 231142 119144 232630 119354
rect 232798 119144 234194 119354
rect 234362 119144 235850 119354
rect 236018 119144 237414 119354
rect 237582 119144 239070 119354
rect 756 856 239180 119144
rect 756 734 790 856
rect 958 734 2446 856
rect 2614 734 4102 856
rect 4270 734 5758 856
rect 5926 734 7414 856
rect 7582 734 9162 856
rect 9330 734 10818 856
rect 10986 734 12474 856
rect 12642 734 14130 856
rect 14298 734 15878 856
rect 16046 734 17534 856
rect 17702 734 19190 856
rect 19358 734 20846 856
rect 21014 734 22594 856
rect 22762 734 24250 856
rect 24418 734 25906 856
rect 26074 734 27562 856
rect 27730 734 29310 856
rect 29478 734 30966 856
rect 31134 734 32622 856
rect 32790 734 34278 856
rect 34446 734 36026 856
rect 36194 734 37682 856
rect 37850 734 39338 856
rect 39506 734 40994 856
rect 41162 734 42742 856
rect 42910 734 44398 856
rect 44566 734 46054 856
rect 46222 734 47710 856
rect 47878 734 49458 856
rect 49626 734 51114 856
rect 51282 734 52770 856
rect 52938 734 54426 856
rect 54594 734 56174 856
rect 56342 734 57830 856
rect 57998 734 59486 856
rect 59654 734 61142 856
rect 61310 734 62890 856
rect 63058 734 64546 856
rect 64714 734 66202 856
rect 66370 734 67858 856
rect 68026 734 69606 856
rect 69774 734 71262 856
rect 71430 734 72918 856
rect 73086 734 74574 856
rect 74742 734 76322 856
rect 76490 734 77978 856
rect 78146 734 79634 856
rect 79802 734 81290 856
rect 81458 734 82946 856
rect 83114 734 84694 856
rect 84862 734 86350 856
rect 86518 734 88006 856
rect 88174 734 89662 856
rect 89830 734 91410 856
rect 91578 734 93066 856
rect 93234 734 94722 856
rect 94890 734 96378 856
rect 96546 734 98126 856
rect 98294 734 99782 856
rect 99950 734 101438 856
rect 101606 734 103094 856
rect 103262 734 104842 856
rect 105010 734 106498 856
rect 106666 734 108154 856
rect 108322 734 109810 856
rect 109978 734 111558 856
rect 111726 734 113214 856
rect 113382 734 114870 856
rect 115038 734 116526 856
rect 116694 734 118274 856
rect 118442 734 119930 856
rect 120098 734 121586 856
rect 121754 734 123242 856
rect 123410 734 124990 856
rect 125158 734 126646 856
rect 126814 734 128302 856
rect 128470 734 129958 856
rect 130126 734 131706 856
rect 131874 734 133362 856
rect 133530 734 135018 856
rect 135186 734 136674 856
rect 136842 734 138422 856
rect 138590 734 140078 856
rect 140246 734 141734 856
rect 141902 734 143390 856
rect 143558 734 145138 856
rect 145306 734 146794 856
rect 146962 734 148450 856
rect 148618 734 150106 856
rect 150274 734 151854 856
rect 152022 734 153510 856
rect 153678 734 155166 856
rect 155334 734 156822 856
rect 156990 734 158570 856
rect 158738 734 160226 856
rect 160394 734 161882 856
rect 162050 734 163538 856
rect 163706 734 165194 856
rect 165362 734 166942 856
rect 167110 734 168598 856
rect 168766 734 170254 856
rect 170422 734 171910 856
rect 172078 734 173658 856
rect 173826 734 175314 856
rect 175482 734 176970 856
rect 177138 734 178626 856
rect 178794 734 180374 856
rect 180542 734 182030 856
rect 182198 734 183686 856
rect 183854 734 185342 856
rect 185510 734 187090 856
rect 187258 734 188746 856
rect 188914 734 190402 856
rect 190570 734 192058 856
rect 192226 734 193806 856
rect 193974 734 195462 856
rect 195630 734 197118 856
rect 197286 734 198774 856
rect 198942 734 200522 856
rect 200690 734 202178 856
rect 202346 734 203834 856
rect 204002 734 205490 856
rect 205658 734 207238 856
rect 207406 734 208894 856
rect 209062 734 210550 856
rect 210718 734 212206 856
rect 212374 734 213954 856
rect 214122 734 215610 856
rect 215778 734 217266 856
rect 217434 734 218922 856
rect 219090 734 220670 856
rect 220838 734 222326 856
rect 222494 734 223982 856
rect 224150 734 225638 856
rect 225806 734 227386 856
rect 227554 734 229042 856
rect 229210 734 230698 856
rect 230866 734 232354 856
rect 232522 734 234102 856
rect 234270 734 235758 856
rect 235926 734 237414 856
rect 237582 734 239070 856
<< metal3 >>
rect 0 117920 800 118040
rect 239200 117512 240000 117632
rect 0 114112 800 114232
rect 239200 112888 240000 113008
rect 0 110440 800 110560
rect 239200 108264 240000 108384
rect 0 106632 800 106752
rect 239200 103640 240000 103760
rect 0 102960 800 103080
rect 0 99152 800 99272
rect 239200 99016 240000 99136
rect 0 95480 800 95600
rect 239200 94392 240000 94512
rect 0 91672 800 91792
rect 239200 89768 240000 89888
rect 0 87864 800 87984
rect 239200 85144 240000 85264
rect 0 84192 800 84312
rect 0 80384 800 80504
rect 239200 80520 240000 80640
rect 0 76712 800 76832
rect 239200 75896 240000 76016
rect 0 72904 800 73024
rect 239200 71272 240000 71392
rect 0 69232 800 69352
rect 239200 66648 240000 66768
rect 0 65424 800 65544
rect 239200 62160 240000 62280
rect 0 61752 800 61872
rect 0 57944 800 58064
rect 239200 57536 240000 57656
rect 0 54136 800 54256
rect 239200 52912 240000 53032
rect 0 50464 800 50584
rect 239200 48288 240000 48408
rect 0 46656 800 46776
rect 239200 43664 240000 43784
rect 0 42984 800 43104
rect 0 39176 800 39296
rect 239200 39040 240000 39160
rect 0 35504 800 35624
rect 239200 34416 240000 34536
rect 0 31696 800 31816
rect 239200 29792 240000 29912
rect 0 27888 800 28008
rect 239200 25168 240000 25288
rect 0 24216 800 24336
rect 0 20408 800 20528
rect 239200 20544 240000 20664
rect 0 16736 800 16856
rect 239200 15920 240000 16040
rect 0 12928 800 13048
rect 239200 11296 240000 11416
rect 0 9256 800 9376
rect 239200 6672 240000 6792
rect 0 5448 800 5568
rect 239200 2184 240000 2304
rect 0 1776 800 1896
<< obsm3 >>
rect 880 117840 239200 118013
rect 800 117712 239200 117840
rect 800 117432 239120 117712
rect 800 114312 239200 117432
rect 880 114032 239200 114312
rect 800 113088 239200 114032
rect 800 112808 239120 113088
rect 800 110640 239200 112808
rect 880 110360 239200 110640
rect 800 108464 239200 110360
rect 800 108184 239120 108464
rect 800 106832 239200 108184
rect 880 106552 239200 106832
rect 800 103840 239200 106552
rect 800 103560 239120 103840
rect 800 103160 239200 103560
rect 880 102880 239200 103160
rect 800 99352 239200 102880
rect 880 99216 239200 99352
rect 880 99072 239120 99216
rect 800 98936 239120 99072
rect 800 95680 239200 98936
rect 880 95400 239200 95680
rect 800 94592 239200 95400
rect 800 94312 239120 94592
rect 800 91872 239200 94312
rect 880 91592 239200 91872
rect 800 89968 239200 91592
rect 800 89688 239120 89968
rect 800 88064 239200 89688
rect 880 87784 239200 88064
rect 800 85344 239200 87784
rect 800 85064 239120 85344
rect 800 84392 239200 85064
rect 880 84112 239200 84392
rect 800 80720 239200 84112
rect 800 80584 239120 80720
rect 880 80440 239120 80584
rect 880 80304 239200 80440
rect 800 76912 239200 80304
rect 880 76632 239200 76912
rect 800 76096 239200 76632
rect 800 75816 239120 76096
rect 800 73104 239200 75816
rect 880 72824 239200 73104
rect 800 71472 239200 72824
rect 800 71192 239120 71472
rect 800 69432 239200 71192
rect 880 69152 239200 69432
rect 800 66848 239200 69152
rect 800 66568 239120 66848
rect 800 65624 239200 66568
rect 880 65344 239200 65624
rect 800 62360 239200 65344
rect 800 62080 239120 62360
rect 800 61952 239200 62080
rect 880 61672 239200 61952
rect 800 58144 239200 61672
rect 880 57864 239200 58144
rect 800 57736 239200 57864
rect 800 57456 239120 57736
rect 800 54336 239200 57456
rect 880 54056 239200 54336
rect 800 53112 239200 54056
rect 800 52832 239120 53112
rect 800 50664 239200 52832
rect 880 50384 239200 50664
rect 800 48488 239200 50384
rect 800 48208 239120 48488
rect 800 46856 239200 48208
rect 880 46576 239200 46856
rect 800 43864 239200 46576
rect 800 43584 239120 43864
rect 800 43184 239200 43584
rect 880 42904 239200 43184
rect 800 39376 239200 42904
rect 880 39240 239200 39376
rect 880 39096 239120 39240
rect 800 38960 239120 39096
rect 800 35704 239200 38960
rect 880 35424 239200 35704
rect 800 34616 239200 35424
rect 800 34336 239120 34616
rect 800 31896 239200 34336
rect 880 31616 239200 31896
rect 800 29992 239200 31616
rect 800 29712 239120 29992
rect 800 28088 239200 29712
rect 880 27808 239200 28088
rect 800 25368 239200 27808
rect 800 25088 239120 25368
rect 800 24416 239200 25088
rect 880 24136 239200 24416
rect 800 20744 239200 24136
rect 800 20608 239120 20744
rect 880 20464 239120 20608
rect 880 20328 239200 20464
rect 800 16936 239200 20328
rect 880 16656 239200 16936
rect 800 16120 239200 16656
rect 800 15840 239120 16120
rect 800 13128 239200 15840
rect 880 12848 239200 13128
rect 800 11496 239200 12848
rect 800 11216 239120 11496
rect 800 9456 239200 11216
rect 880 9176 239200 9456
rect 800 6872 239200 9176
rect 800 6592 239120 6872
rect 800 5648 239200 6592
rect 880 5368 239200 5648
rect 800 2384 239200 5368
rect 800 2104 239120 2384
rect 800 1976 239200 2104
rect 880 1803 239200 1976
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
rect 188528 2128 188848 117552
rect 203888 2128 204208 117552
rect 219248 2128 219568 117552
rect 234608 2128 234928 117552
<< obsm4 >>
rect 58203 11731 65568 109717
rect 66048 11731 80928 109717
rect 81408 11731 96288 109717
rect 96768 11731 111648 109717
rect 112128 11731 127008 109717
rect 127488 11731 142368 109717
rect 142848 11731 157728 109717
rect 158208 11731 173088 109717
rect 173568 11731 188448 109717
rect 188928 11731 203808 109717
rect 204288 11731 213749 109717
<< labels >>
rlabel metal2 s 10414 119200 10470 120000 6 addrA0[0]
port 1 nsew signal output
rlabel metal2 s 11978 119200 12034 120000 6 addrA0[1]
port 2 nsew signal output
rlabel metal2 s 13634 119200 13690 120000 6 addrA0[2]
port 3 nsew signal output
rlabel metal2 s 15198 119200 15254 120000 6 addrA0[3]
port 4 nsew signal output
rlabel metal2 s 16854 119200 16910 120000 6 addrA0[4]
port 5 nsew signal output
rlabel metal2 s 18418 119200 18474 120000 6 addrA0[5]
port 6 nsew signal output
rlabel metal2 s 20074 119200 20130 120000 6 addrA0[6]
port 7 nsew signal output
rlabel metal2 s 21638 119200 21694 120000 6 addrA0[7]
port 8 nsew signal output
rlabel metal2 s 23294 119200 23350 120000 6 addrA1[0]
port 9 nsew signal output
rlabel metal2 s 24858 119200 24914 120000 6 addrA1[1]
port 10 nsew signal output
rlabel metal2 s 26514 119200 26570 120000 6 addrA1[2]
port 11 nsew signal output
rlabel metal2 s 28078 119200 28134 120000 6 addrA1[3]
port 12 nsew signal output
rlabel metal2 s 29734 119200 29790 120000 6 addrA1[4]
port 13 nsew signal output
rlabel metal2 s 31298 119200 31354 120000 6 addrA1[5]
port 14 nsew signal output
rlabel metal2 s 32954 119200 33010 120000 6 addrA1[6]
port 15 nsew signal output
rlabel metal2 s 34518 119200 34574 120000 6 addrA1[7]
port 16 nsew signal output
rlabel metal2 s 94134 119200 94190 120000 6 addrB0[0]
port 17 nsew signal output
rlabel metal2 s 95790 119200 95846 120000 6 addrB0[1]
port 18 nsew signal output
rlabel metal2 s 97354 119200 97410 120000 6 addrB0[2]
port 19 nsew signal output
rlabel metal2 s 99010 119200 99066 120000 6 addrB0[3]
port 20 nsew signal output
rlabel metal2 s 100574 119200 100630 120000 6 addrB0[4]
port 21 nsew signal output
rlabel metal2 s 102230 119200 102286 120000 6 addrB0[5]
port 22 nsew signal output
rlabel metal2 s 103794 119200 103850 120000 6 addrB0[6]
port 23 nsew signal output
rlabel metal2 s 105450 119200 105506 120000 6 addrB0[7]
port 24 nsew signal output
rlabel metal2 s 107014 119200 107070 120000 6 addrB0[8]
port 25 nsew signal output
rlabel metal2 s 108670 119200 108726 120000 6 addrB1[0]
port 26 nsew signal output
rlabel metal2 s 110234 119200 110290 120000 6 addrB1[1]
port 27 nsew signal output
rlabel metal2 s 111890 119200 111946 120000 6 addrB1[2]
port 28 nsew signal output
rlabel metal2 s 113454 119200 113510 120000 6 addrB1[3]
port 29 nsew signal output
rlabel metal2 s 115110 119200 115166 120000 6 addrB1[4]
port 30 nsew signal output
rlabel metal2 s 116674 119200 116730 120000 6 addrB1[5]
port 31 nsew signal output
rlabel metal2 s 118330 119200 118386 120000 6 addrB1[6]
port 32 nsew signal output
rlabel metal2 s 119894 119200 119950 120000 6 addrB1[7]
port 33 nsew signal output
rlabel metal2 s 121550 119200 121606 120000 6 addrB1[8]
port 34 nsew signal output
rlabel metal2 s 7194 119200 7250 120000 6 csbA0
port 35 nsew signal output
rlabel metal2 s 8758 119200 8814 120000 6 csbA1
port 36 nsew signal output
rlabel metal2 s 754 119200 810 120000 6 csbB0
port 37 nsew signal output
rlabel metal2 s 2318 119200 2374 120000 6 csbB1
port 38 nsew signal output
rlabel metal2 s 36174 119200 36230 120000 6 dinA0[0]
port 39 nsew signal output
rlabel metal2 s 52274 119200 52330 120000 6 dinA0[10]
port 40 nsew signal output
rlabel metal2 s 53838 119200 53894 120000 6 dinA0[11]
port 41 nsew signal output
rlabel metal2 s 55494 119200 55550 120000 6 dinA0[12]
port 42 nsew signal output
rlabel metal2 s 57058 119200 57114 120000 6 dinA0[13]
port 43 nsew signal output
rlabel metal2 s 58714 119200 58770 120000 6 dinA0[14]
port 44 nsew signal output
rlabel metal2 s 60278 119200 60334 120000 6 dinA0[15]
port 45 nsew signal output
rlabel metal2 s 61934 119200 61990 120000 6 dinA0[16]
port 46 nsew signal output
rlabel metal2 s 63498 119200 63554 120000 6 dinA0[17]
port 47 nsew signal output
rlabel metal2 s 65154 119200 65210 120000 6 dinA0[18]
port 48 nsew signal output
rlabel metal2 s 66718 119200 66774 120000 6 dinA0[19]
port 49 nsew signal output
rlabel metal2 s 37738 119200 37794 120000 6 dinA0[1]
port 50 nsew signal output
rlabel metal2 s 68374 119200 68430 120000 6 dinA0[20]
port 51 nsew signal output
rlabel metal2 s 69938 119200 69994 120000 6 dinA0[21]
port 52 nsew signal output
rlabel metal2 s 71594 119200 71650 120000 6 dinA0[22]
port 53 nsew signal output
rlabel metal2 s 73158 119200 73214 120000 6 dinA0[23]
port 54 nsew signal output
rlabel metal2 s 74814 119200 74870 120000 6 dinA0[24]
port 55 nsew signal output
rlabel metal2 s 76378 119200 76434 120000 6 dinA0[25]
port 56 nsew signal output
rlabel metal2 s 78034 119200 78090 120000 6 dinA0[26]
port 57 nsew signal output
rlabel metal2 s 79598 119200 79654 120000 6 dinA0[27]
port 58 nsew signal output
rlabel metal2 s 81254 119200 81310 120000 6 dinA0[28]
port 59 nsew signal output
rlabel metal2 s 82910 119200 82966 120000 6 dinA0[29]
port 60 nsew signal output
rlabel metal2 s 39394 119200 39450 120000 6 dinA0[2]
port 61 nsew signal output
rlabel metal2 s 84474 119200 84530 120000 6 dinA0[30]
port 62 nsew signal output
rlabel metal2 s 86130 119200 86186 120000 6 dinA0[31]
port 63 nsew signal output
rlabel metal2 s 40958 119200 41014 120000 6 dinA0[3]
port 64 nsew signal output
rlabel metal2 s 42614 119200 42670 120000 6 dinA0[4]
port 65 nsew signal output
rlabel metal2 s 44178 119200 44234 120000 6 dinA0[5]
port 66 nsew signal output
rlabel metal2 s 45834 119200 45890 120000 6 dinA0[6]
port 67 nsew signal output
rlabel metal2 s 47398 119200 47454 120000 6 dinA0[7]
port 68 nsew signal output
rlabel metal2 s 49054 119200 49110 120000 6 dinA0[8]
port 69 nsew signal output
rlabel metal2 s 50618 119200 50674 120000 6 dinA0[9]
port 70 nsew signal output
rlabel metal2 s 123114 119200 123170 120000 6 dinB0[0]
port 71 nsew signal output
rlabel metal2 s 139214 119200 139270 120000 6 dinB0[10]
port 72 nsew signal output
rlabel metal2 s 140870 119200 140926 120000 6 dinB0[11]
port 73 nsew signal output
rlabel metal2 s 142434 119200 142490 120000 6 dinB0[12]
port 74 nsew signal output
rlabel metal2 s 144090 119200 144146 120000 6 dinB0[13]
port 75 nsew signal output
rlabel metal2 s 145654 119200 145710 120000 6 dinB0[14]
port 76 nsew signal output
rlabel metal2 s 147310 119200 147366 120000 6 dinB0[15]
port 77 nsew signal output
rlabel metal2 s 148874 119200 148930 120000 6 dinB0[16]
port 78 nsew signal output
rlabel metal2 s 150530 119200 150586 120000 6 dinB0[17]
port 79 nsew signal output
rlabel metal2 s 152094 119200 152150 120000 6 dinB0[18]
port 80 nsew signal output
rlabel metal2 s 153750 119200 153806 120000 6 dinB0[19]
port 81 nsew signal output
rlabel metal2 s 124770 119200 124826 120000 6 dinB0[1]
port 82 nsew signal output
rlabel metal2 s 155314 119200 155370 120000 6 dinB0[20]
port 83 nsew signal output
rlabel metal2 s 156970 119200 157026 120000 6 dinB0[21]
port 84 nsew signal output
rlabel metal2 s 158534 119200 158590 120000 6 dinB0[22]
port 85 nsew signal output
rlabel metal2 s 160190 119200 160246 120000 6 dinB0[23]
port 86 nsew signal output
rlabel metal2 s 161846 119200 161902 120000 6 dinB0[24]
port 87 nsew signal output
rlabel metal2 s 163410 119200 163466 120000 6 dinB0[25]
port 88 nsew signal output
rlabel metal2 s 165066 119200 165122 120000 6 dinB0[26]
port 89 nsew signal output
rlabel metal2 s 166630 119200 166686 120000 6 dinB0[27]
port 90 nsew signal output
rlabel metal2 s 168286 119200 168342 120000 6 dinB0[28]
port 91 nsew signal output
rlabel metal2 s 169850 119200 169906 120000 6 dinB0[29]
port 92 nsew signal output
rlabel metal2 s 126334 119200 126390 120000 6 dinB0[2]
port 93 nsew signal output
rlabel metal2 s 171506 119200 171562 120000 6 dinB0[30]
port 94 nsew signal output
rlabel metal2 s 173070 119200 173126 120000 6 dinB0[31]
port 95 nsew signal output
rlabel metal2 s 127990 119200 128046 120000 6 dinB0[3]
port 96 nsew signal output
rlabel metal2 s 129554 119200 129610 120000 6 dinB0[4]
port 97 nsew signal output
rlabel metal2 s 131210 119200 131266 120000 6 dinB0[5]
port 98 nsew signal output
rlabel metal2 s 132774 119200 132830 120000 6 dinB0[6]
port 99 nsew signal output
rlabel metal2 s 134430 119200 134486 120000 6 dinB0[7]
port 100 nsew signal output
rlabel metal2 s 135994 119200 136050 120000 6 dinB0[8]
port 101 nsew signal output
rlabel metal2 s 137650 119200 137706 120000 6 dinB0[9]
port 102 nsew signal output
rlabel metal2 s 182730 119200 182786 120000 6 sram12_dout0[0]
port 103 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 sram12_dout0[10]
port 104 nsew signal input
rlabel metal3 s 239200 57536 240000 57656 6 sram12_dout0[11]
port 105 nsew signal input
rlabel metal2 s 200486 119200 200542 120000 6 sram12_dout0[12]
port 106 nsew signal input
rlabel metal2 s 207294 0 207350 800 6 sram12_dout0[13]
port 107 nsew signal input
rlabel metal2 s 206926 119200 206982 120000 6 sram12_dout0[14]
port 108 nsew signal input
rlabel metal2 s 212262 0 212318 800 6 sram12_dout0[15]
port 109 nsew signal input
rlabel metal2 s 208490 119200 208546 120000 6 sram12_dout0[16]
port 110 nsew signal input
rlabel metal2 s 210146 119200 210202 120000 6 sram12_dout0[17]
port 111 nsew signal input
rlabel metal3 s 239200 75896 240000 76016 6 sram12_dout0[18]
port 112 nsew signal input
rlabel metal2 s 222382 0 222438 800 6 sram12_dout0[19]
port 113 nsew signal input
rlabel metal2 s 180430 0 180486 800 6 sram12_dout0[1]
port 114 nsew signal input
rlabel metal2 s 214930 119200 214986 120000 6 sram12_dout0[20]
port 115 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 sram12_dout0[21]
port 116 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 sram12_dout0[22]
port 117 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 sram12_dout0[23]
port 118 nsew signal input
rlabel metal2 s 230754 0 230810 800 6 sram12_dout0[24]
port 119 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 sram12_dout0[25]
port 120 nsew signal input
rlabel metal2 s 227810 119200 227866 120000 6 sram12_dout0[26]
port 121 nsew signal input
rlabel metal2 s 231030 119200 231086 120000 6 sram12_dout0[27]
port 122 nsew signal input
rlabel metal2 s 234158 0 234214 800 6 sram12_dout0[28]
port 123 nsew signal input
rlabel metal2 s 237470 0 237526 800 6 sram12_dout0[29]
port 124 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 sram12_dout0[2]
port 125 nsew signal input
rlabel metal2 s 237470 119200 237526 120000 6 sram12_dout0[30]
port 126 nsew signal input
rlabel metal3 s 239200 117512 240000 117632 6 sram12_dout0[31]
port 127 nsew signal input
rlabel metal2 s 187606 119200 187662 120000 6 sram12_dout0[3]
port 128 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 sram12_dout0[4]
port 129 nsew signal input
rlabel metal2 s 192114 0 192170 800 6 sram12_dout0[5]
port 130 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 sram12_dout0[6]
port 131 nsew signal input
rlabel metal2 s 197174 0 197230 800 6 sram12_dout0[7]
port 132 nsew signal input
rlabel metal2 s 194046 119200 194102 120000 6 sram12_dout0[8]
port 133 nsew signal input
rlabel metal2 s 195610 119200 195666 120000 6 sram12_dout0[9]
port 134 nsew signal input
rlabel metal2 s 184386 119200 184442 120000 6 sram12_dout1[0]
port 135 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 sram12_dout1[10]
port 136 nsew signal input
rlabel metal2 s 198830 119200 198886 120000 6 sram12_dout1[11]
port 137 nsew signal input
rlabel metal2 s 202050 119200 202106 120000 6 sram12_dout1[12]
port 138 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 sram12_dout1[13]
port 139 nsew signal input
rlabel metal3 s 239200 62160 240000 62280 6 sram12_dout1[14]
port 140 nsew signal input
rlabel metal3 s 239200 66648 240000 66768 6 sram12_dout1[15]
port 141 nsew signal input
rlabel metal2 s 215666 0 215722 800 6 sram12_dout1[16]
port 142 nsew signal input
rlabel metal2 s 217322 0 217378 800 6 sram12_dout1[17]
port 143 nsew signal input
rlabel metal2 s 213366 119200 213422 120000 6 sram12_dout1[18]
port 144 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 sram12_dout1[19]
port 145 nsew signal input
rlabel metal3 s 239200 6672 240000 6792 6 sram12_dout1[1]
port 146 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 sram12_dout1[20]
port 147 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 sram12_dout1[21]
port 148 nsew signal input
rlabel metal2 s 221370 119200 221426 120000 6 sram12_dout1[22]
port 149 nsew signal input
rlabel metal2 s 223026 119200 223082 120000 6 sram12_dout1[23]
port 150 nsew signal input
rlabel metal2 s 224590 119200 224646 120000 6 sram12_dout1[24]
port 151 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 sram12_dout1[25]
port 152 nsew signal input
rlabel metal3 s 239200 103640 240000 103760 6 sram12_dout1[26]
port 153 nsew signal input
rlabel metal2 s 232686 119200 232742 120000 6 sram12_dout1[27]
port 154 nsew signal input
rlabel metal2 s 235814 0 235870 800 6 sram12_dout1[28]
port 155 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 sram12_dout1[29]
port 156 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 sram12_dout1[2]
port 157 nsew signal input
rlabel metal3 s 239200 112888 240000 113008 6 sram12_dout1[30]
port 158 nsew signal input
rlabel metal2 s 239126 119200 239182 120000 6 sram12_dout1[31]
port 159 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 sram12_dout1[3]
port 160 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 sram12_dout1[4]
port 161 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 sram12_dout1[5]
port 162 nsew signal input
rlabel metal2 s 192390 119200 192446 120000 6 sram12_dout1[6]
port 163 nsew signal input
rlabel metal3 s 239200 34416 240000 34536 6 sram12_dout1[7]
port 164 nsew signal input
rlabel metal3 s 239200 39040 240000 39160 6 sram12_dout1[8]
port 165 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 sram12_dout1[9]
port 166 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 sram1_dout0[0]
port 167 nsew signal input
rlabel metal2 s 197266 119200 197322 120000 6 sram1_dout0[10]
port 168 nsew signal input
rlabel metal3 s 239200 48288 240000 48408 6 sram1_dout0[11]
port 169 nsew signal input
rlabel metal2 s 203890 0 203946 800 6 sram1_dout0[12]
port 170 nsew signal input
rlabel metal2 s 203706 119200 203762 120000 6 sram1_dout0[13]
port 171 nsew signal input
rlabel metal2 s 205270 119200 205326 120000 6 sram1_dout0[14]
port 172 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 sram1_dout0[15]
port 173 nsew signal input
rlabel metal3 s 239200 71272 240000 71392 6 sram1_dout0[16]
port 174 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 sram1_dout0[17]
port 175 nsew signal input
rlabel metal2 s 218978 0 219034 800 6 sram1_dout0[18]
port 176 nsew signal input
rlabel metal2 s 220726 0 220782 800 6 sram1_dout0[19]
port 177 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 sram1_dout0[1]
port 178 nsew signal input
rlabel metal2 s 224038 0 224094 800 6 sram1_dout0[20]
port 179 nsew signal input
rlabel metal3 s 239200 85144 240000 85264 6 sram1_dout0[21]
port 180 nsew signal input
rlabel metal2 s 218150 119200 218206 120000 6 sram1_dout0[22]
port 181 nsew signal input
rlabel metal2 s 227442 0 227498 800 6 sram1_dout0[23]
port 182 nsew signal input
rlabel metal2 s 229098 0 229154 800 6 sram1_dout0[24]
port 183 nsew signal input
rlabel metal3 s 239200 89768 240000 89888 6 sram1_dout0[25]
port 184 nsew signal input
rlabel metal2 s 226246 119200 226302 120000 6 sram1_dout0[26]
port 185 nsew signal input
rlabel metal2 s 229466 119200 229522 120000 6 sram1_dout0[27]
port 186 nsew signal input
rlabel metal2 s 232410 0 232466 800 6 sram1_dout0[28]
port 187 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 sram1_dout0[29]
port 188 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 sram1_dout0[2]
port 189 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 sram1_dout0[30]
port 190 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 sram1_dout0[31]
port 191 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 sram1_dout0[3]
port 192 nsew signal input
rlabel metal2 s 189170 119200 189226 120000 6 sram1_dout0[4]
port 193 nsew signal input
rlabel metal2 s 190826 119200 190882 120000 6 sram1_dout0[5]
port 194 nsew signal input
rlabel metal3 s 239200 25168 240000 25288 6 sram1_dout0[6]
port 195 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 sram1_dout0[7]
port 196 nsew signal input
rlabel metal2 s 198830 0 198886 800 6 sram1_dout0[8]
port 197 nsew signal input
rlabel metal2 s 200578 0 200634 800 6 sram1_dout0[9]
port 198 nsew signal input
rlabel metal2 s 181166 119200 181222 120000 6 sram1_dout1[0]
port 199 nsew signal input
rlabel metal3 s 0 35504 800 35624 6 sram1_dout1[10]
port 200 nsew signal input
rlabel metal3 s 239200 52912 240000 53032 6 sram1_dout1[11]
port 201 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 sram1_dout1[12]
port 202 nsew signal input
rlabel metal2 s 205546 0 205602 800 6 sram1_dout1[13]
port 203 nsew signal input
rlabel metal2 s 208950 0 209006 800 6 sram1_dout1[14]
port 204 nsew signal input
rlabel metal2 s 210606 0 210662 800 6 sram1_dout1[15]
port 205 nsew signal input
rlabel metal2 s 214010 0 214066 800 6 sram1_dout1[16]
port 206 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 sram1_dout1[17]
port 207 nsew signal input
rlabel metal2 s 211710 119200 211766 120000 6 sram1_dout1[18]
port 208 nsew signal input
rlabel metal3 s 0 65424 800 65544 6 sram1_dout1[19]
port 209 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 sram1_dout1[1]
port 210 nsew signal input
rlabel metal3 s 239200 80520 240000 80640 6 sram1_dout1[20]
port 211 nsew signal input
rlabel metal2 s 216586 119200 216642 120000 6 sram1_dout1[21]
port 212 nsew signal input
rlabel metal2 s 219806 119200 219862 120000 6 sram1_dout1[22]
port 213 nsew signal input
rlabel metal3 s 0 84192 800 84312 6 sram1_dout1[23]
port 214 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 sram1_dout1[24]
port 215 nsew signal input
rlabel metal3 s 239200 94392 240000 94512 6 sram1_dout1[25]
port 216 nsew signal input
rlabel metal3 s 239200 99016 240000 99136 6 sram1_dout1[26]
port 217 nsew signal input
rlabel metal3 s 239200 108264 240000 108384 6 sram1_dout1[27]
port 218 nsew signal input
rlabel metal2 s 234250 119200 234306 120000 6 sram1_dout1[28]
port 219 nsew signal input
rlabel metal2 s 235906 119200 235962 120000 6 sram1_dout1[29]
port 220 nsew signal input
rlabel metal2 s 185950 119200 186006 120000 6 sram1_dout1[2]
port 221 nsew signal input
rlabel metal2 s 239126 0 239182 800 6 sram1_dout1[30]
port 222 nsew signal input
rlabel metal3 s 0 117920 800 118040 6 sram1_dout1[31]
port 223 nsew signal input
rlabel metal3 s 239200 15920 240000 16040 6 sram1_dout1[3]
port 224 nsew signal input
rlabel metal3 s 239200 20544 240000 20664 6 sram1_dout1[4]
port 225 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 sram1_dout1[5]
port 226 nsew signal input
rlabel metal3 s 239200 29792 240000 29912 6 sram1_dout1[6]
port 227 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 sram1_dout1[7]
port 228 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 sram1_dout1[8]
port 229 nsew signal input
rlabel metal3 s 239200 43664 240000 43784 6 sram1_dout1[9]
port 230 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 user_clock2
port 231 nsew signal input
rlabel metal3 s 239200 2184 240000 2304 6 user_irq[0]
port 232 nsew signal output
rlabel metal3 s 239200 11296 240000 11416 6 user_irq[1]
port 233 nsew signal output
rlabel metal2 s 185398 0 185454 800 6 user_irq[2]
port 234 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 235 nsew power input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 235 nsew power input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 235 nsew power input
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 235 nsew power input
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 235 nsew power input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 235 nsew power input
rlabel metal4 s 188528 2128 188848 117552 6 vccd1
port 235 nsew power input
rlabel metal4 s 219248 2128 219568 117552 6 vccd1
port 235 nsew power input
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 236 nsew ground input
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 236 nsew ground input
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 236 nsew ground input
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 236 nsew ground input
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 236 nsew ground input
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 236 nsew ground input
rlabel metal4 s 203888 2128 204208 117552 6 vssd1
port 236 nsew ground input
rlabel metal4 s 234608 2128 234928 117552 6 vssd1
port 236 nsew ground input
rlabel metal2 s 846 0 902 800 6 wb_clk_i
port 237 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wb_rst_i
port 238 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_ack_o
port 239 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[0]
port 240 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 wbs_adr_i[10]
port 241 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 wbs_adr_i[11]
port 242 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 wbs_adr_i[12]
port 243 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 wbs_adr_i[13]
port 244 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 wbs_adr_i[14]
port 245 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 wbs_adr_i[15]
port 246 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 wbs_adr_i[16]
port 247 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 wbs_adr_i[17]
port 248 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 wbs_adr_i[18]
port 249 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 wbs_adr_i[19]
port 250 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[1]
port 251 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 wbs_adr_i[20]
port 252 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 wbs_adr_i[21]
port 253 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 wbs_adr_i[22]
port 254 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 wbs_adr_i[23]
port 255 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 wbs_adr_i[24]
port 256 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 wbs_adr_i[25]
port 257 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 wbs_adr_i[26]
port 258 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 wbs_adr_i[27]
port 259 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 wbs_adr_i[28]
port 260 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 wbs_adr_i[29]
port 261 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_adr_i[2]
port 262 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 wbs_adr_i[30]
port 263 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 wbs_adr_i[31]
port 264 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[3]
port 265 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_adr_i[4]
port 266 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_adr_i[5]
port 267 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 wbs_adr_i[6]
port 268 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 wbs_adr_i[7]
port 269 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 wbs_adr_i[8]
port 270 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 wbs_adr_i[9]
port 271 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_cyc_i
port 272 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_i[0]
port 273 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 wbs_dat_i[10]
port 274 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 wbs_dat_i[11]
port 275 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 wbs_dat_i[12]
port 276 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 wbs_dat_i[13]
port 277 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 wbs_dat_i[14]
port 278 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 wbs_dat_i[15]
port 279 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 wbs_dat_i[16]
port 280 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 wbs_dat_i[17]
port 281 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 wbs_dat_i[18]
port 282 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 wbs_dat_i[19]
port 283 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[1]
port 284 nsew signal input
rlabel metal2 s 119986 0 120042 800 6 wbs_dat_i[20]
port 285 nsew signal input
rlabel metal2 s 125046 0 125102 800 6 wbs_dat_i[21]
port 286 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 wbs_dat_i[22]
port 287 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 wbs_dat_i[23]
port 288 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 wbs_dat_i[24]
port 289 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 wbs_dat_i[25]
port 290 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 wbs_dat_i[26]
port 291 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 wbs_dat_i[27]
port 292 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 wbs_dat_i[28]
port 293 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 wbs_dat_i[29]
port 294 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_i[2]
port 295 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 wbs_dat_i[30]
port 296 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 wbs_dat_i[31]
port 297 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[3]
port 298 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_i[4]
port 299 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_dat_i[5]
port 300 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 wbs_dat_i[6]
port 301 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 wbs_dat_i[7]
port 302 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_i[8]
port 303 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 wbs_dat_i[9]
port 304 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[0]
port 305 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 wbs_dat_o[10]
port 306 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 wbs_dat_o[11]
port 307 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 wbs_dat_o[12]
port 308 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 wbs_dat_o[13]
port 309 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 wbs_dat_o[14]
port 310 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 wbs_dat_o[15]
port 311 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 wbs_dat_o[16]
port 312 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 wbs_dat_o[17]
port 313 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 wbs_dat_o[18]
port 314 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 wbs_dat_o[19]
port 315 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[1]
port 316 nsew signal output
rlabel metal2 s 121642 0 121698 800 6 wbs_dat_o[20]
port 317 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 wbs_dat_o[21]
port 318 nsew signal output
rlabel metal2 s 131762 0 131818 800 6 wbs_dat_o[22]
port 319 nsew signal output
rlabel metal2 s 136730 0 136786 800 6 wbs_dat_o[23]
port 320 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 wbs_dat_o[24]
port 321 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 wbs_dat_o[25]
port 322 nsew signal output
rlabel metal2 s 151910 0 151966 800 6 wbs_dat_o[26]
port 323 nsew signal output
rlabel metal2 s 156878 0 156934 800 6 wbs_dat_o[27]
port 324 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 wbs_dat_o[28]
port 325 nsew signal output
rlabel metal2 s 166998 0 167054 800 6 wbs_dat_o[29]
port 326 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[2]
port 327 nsew signal output
rlabel metal2 s 171966 0 172022 800 6 wbs_dat_o[30]
port 328 nsew signal output
rlabel metal2 s 177026 0 177082 800 6 wbs_dat_o[31]
port 329 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_o[3]
port 330 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_o[4]
port 331 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_o[5]
port 332 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_o[6]
port 333 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 wbs_dat_o[7]
port 334 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 wbs_dat_o[8]
port 335 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 wbs_dat_o[9]
port 336 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_sel_i[0]
port 337 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_sel_i[1]
port 338 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_sel_i[2]
port 339 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_sel_i[3]
port 340 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_stb_i
port 341 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_we_i
port 342 nsew signal input
rlabel metal2 s 3974 119200 4030 120000 6 webA
port 343 nsew signal output
rlabel metal2 s 5538 119200 5594 120000 6 webB
port 344 nsew signal output
rlabel metal2 s 87694 119200 87750 120000 6 wmaskA[0]
port 345 nsew signal output
rlabel metal2 s 89350 119200 89406 120000 6 wmaskA[1]
port 346 nsew signal output
rlabel metal2 s 90914 119200 90970 120000 6 wmaskA[2]
port 347 nsew signal output
rlabel metal2 s 92570 119200 92626 120000 6 wmaskA[3]
port 348 nsew signal output
rlabel metal2 s 174726 119200 174782 120000 6 wmaskB[0]
port 349 nsew signal output
rlabel metal2 s 176290 119200 176346 120000 6 wmaskB[1]
port 350 nsew signal output
rlabel metal2 s 177946 119200 178002 120000 6 wmaskB[2]
port 351 nsew signal output
rlabel metal2 s 179510 119200 179566 120000 6 wmaskB[3]
port 352 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 240000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 27853394
string GDS_FILE /home/re19/Caravel/temporal_runtime_monitor/openlane/user_project/runs/user_project/results/finishing/user_project.magic.gds
string GDS_START 1676704
<< end >>

