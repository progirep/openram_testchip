magic
tech sky130A
magscale 1 2
timestamp 1649963323
<< obsli1 >>
rect 1104 2159 74888 80529
<< obsm1 >>
rect 14 8 75978 81048
<< metal2 >>
rect 294 82000 350 82800
rect 938 82000 994 82800
rect 1674 82000 1730 82800
rect 2318 82000 2374 82800
rect 3054 82000 3110 82800
rect 3698 82000 3754 82800
rect 4434 82000 4490 82800
rect 5078 82000 5134 82800
rect 5814 82000 5870 82800
rect 6458 82000 6514 82800
rect 7194 82000 7250 82800
rect 7838 82000 7894 82800
rect 8574 82000 8630 82800
rect 9218 82000 9274 82800
rect 9954 82000 10010 82800
rect 10598 82000 10654 82800
rect 11334 82000 11390 82800
rect 11978 82000 12034 82800
rect 12714 82000 12770 82800
rect 13358 82000 13414 82800
rect 14094 82000 14150 82800
rect 14738 82000 14794 82800
rect 15474 82000 15530 82800
rect 16118 82000 16174 82800
rect 16854 82000 16910 82800
rect 17498 82000 17554 82800
rect 18234 82000 18290 82800
rect 18878 82000 18934 82800
rect 19614 82000 19670 82800
rect 20258 82000 20314 82800
rect 20994 82000 21050 82800
rect 21638 82000 21694 82800
rect 22374 82000 22430 82800
rect 23018 82000 23074 82800
rect 23754 82000 23810 82800
rect 24398 82000 24454 82800
rect 25134 82000 25190 82800
rect 25778 82000 25834 82800
rect 26514 82000 26570 82800
rect 27158 82000 27214 82800
rect 27894 82000 27950 82800
rect 28538 82000 28594 82800
rect 29274 82000 29330 82800
rect 29918 82000 29974 82800
rect 30654 82000 30710 82800
rect 31298 82000 31354 82800
rect 32034 82000 32090 82800
rect 32678 82000 32734 82800
rect 33414 82000 33470 82800
rect 34058 82000 34114 82800
rect 34794 82000 34850 82800
rect 35438 82000 35494 82800
rect 36174 82000 36230 82800
rect 36818 82000 36874 82800
rect 37554 82000 37610 82800
rect 38290 82000 38346 82800
rect 38934 82000 38990 82800
rect 39670 82000 39726 82800
rect 40314 82000 40370 82800
rect 41050 82000 41106 82800
rect 41694 82000 41750 82800
rect 42430 82000 42486 82800
rect 43074 82000 43130 82800
rect 43810 82000 43866 82800
rect 44454 82000 44510 82800
rect 45190 82000 45246 82800
rect 45834 82000 45890 82800
rect 46570 82000 46626 82800
rect 47214 82000 47270 82800
rect 47950 82000 48006 82800
rect 48594 82000 48650 82800
rect 49330 82000 49386 82800
rect 49974 82000 50030 82800
rect 50710 82000 50766 82800
rect 51354 82000 51410 82800
rect 52090 82000 52146 82800
rect 52734 82000 52790 82800
rect 53470 82000 53526 82800
rect 54114 82000 54170 82800
rect 54850 82000 54906 82800
rect 55494 82000 55550 82800
rect 56230 82000 56286 82800
rect 56874 82000 56930 82800
rect 57610 82000 57666 82800
rect 58254 82000 58310 82800
rect 58990 82000 59046 82800
rect 59634 82000 59690 82800
rect 60370 82000 60426 82800
rect 61014 82000 61070 82800
rect 61750 82000 61806 82800
rect 62394 82000 62450 82800
rect 63130 82000 63186 82800
rect 63774 82000 63830 82800
rect 64510 82000 64566 82800
rect 65154 82000 65210 82800
rect 65890 82000 65946 82800
rect 66534 82000 66590 82800
rect 67270 82000 67326 82800
rect 67914 82000 67970 82800
rect 68650 82000 68706 82800
rect 69294 82000 69350 82800
rect 70030 82000 70086 82800
rect 70674 82000 70730 82800
rect 71410 82000 71466 82800
rect 72054 82000 72110 82800
rect 72790 82000 72846 82800
rect 73434 82000 73490 82800
rect 74170 82000 74226 82800
rect 74814 82000 74870 82800
rect 75550 82000 75606 82800
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11610 0 11666 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22650 0 22706 800
rect 23018 0 23074 800
rect 23478 0 23534 800
rect 23846 0 23902 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25502 0 25558 800
rect 25870 0 25926 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27894 0 27950 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 30010 0 30066 800
rect 30378 0 30434 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 32034 0 32090 800
rect 32402 0 32458 800
rect 32862 0 32918 800
rect 33230 0 33286 800
rect 33690 0 33746 800
rect 34058 0 34114 800
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35254 0 35310 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37370 0 37426 800
rect 37738 0 37794 800
rect 38198 0 38254 800
rect 38566 0 38622 800
rect 38934 0 38990 800
rect 39394 0 39450 800
rect 39762 0 39818 800
rect 40222 0 40278 800
rect 40590 0 40646 800
rect 41050 0 41106 800
rect 41418 0 41474 800
rect 41786 0 41842 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 43074 0 43130 800
rect 43442 0 43498 800
rect 43902 0 43958 800
rect 44270 0 44326 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45466 0 45522 800
rect 45926 0 45982 800
rect 46294 0 46350 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48410 0 48466 800
rect 48778 0 48834 800
rect 49146 0 49202 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50434 0 50490 800
rect 50802 0 50858 800
rect 51262 0 51318 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53286 0 53342 800
rect 53654 0 53710 800
rect 54114 0 54170 800
rect 54482 0 54538 800
rect 54942 0 54998 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56506 0 56562 800
rect 56966 0 57022 800
rect 57334 0 57390 800
rect 57794 0 57850 800
rect 58162 0 58218 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60646 0 60702 800
rect 61014 0 61070 800
rect 61474 0 61530 800
rect 61842 0 61898 800
rect 62302 0 62358 800
rect 62670 0 62726 800
rect 63038 0 63094 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64326 0 64382 800
rect 64694 0 64750 800
rect 65154 0 65210 800
rect 65522 0 65578 800
rect 65890 0 65946 800
rect 66350 0 66406 800
rect 66718 0 66774 800
rect 67178 0 67234 800
rect 67546 0 67602 800
rect 68006 0 68062 800
rect 68374 0 68430 800
rect 68834 0 68890 800
rect 69202 0 69258 800
rect 69570 0 69626 800
rect 70030 0 70086 800
rect 70398 0 70454 800
rect 70858 0 70914 800
rect 71226 0 71282 800
rect 71686 0 71742 800
rect 72054 0 72110 800
rect 72514 0 72570 800
rect 72882 0 72938 800
rect 73250 0 73306 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75366 0 75422 800
rect 75734 0 75790 800
<< obsm2 >>
rect 20 81944 238 82090
rect 406 81944 882 82090
rect 1050 81944 1618 82090
rect 1786 81944 2262 82090
rect 2430 81944 2998 82090
rect 3166 81944 3642 82090
rect 3810 81944 4378 82090
rect 4546 81944 5022 82090
rect 5190 81944 5758 82090
rect 5926 81944 6402 82090
rect 6570 81944 7138 82090
rect 7306 81944 7782 82090
rect 7950 81944 8518 82090
rect 8686 81944 9162 82090
rect 9330 81944 9898 82090
rect 10066 81944 10542 82090
rect 10710 81944 11278 82090
rect 11446 81944 11922 82090
rect 12090 81944 12658 82090
rect 12826 81944 13302 82090
rect 13470 81944 14038 82090
rect 14206 81944 14682 82090
rect 14850 81944 15418 82090
rect 15586 81944 16062 82090
rect 16230 81944 16798 82090
rect 16966 81944 17442 82090
rect 17610 81944 18178 82090
rect 18346 81944 18822 82090
rect 18990 81944 19558 82090
rect 19726 81944 20202 82090
rect 20370 81944 20938 82090
rect 21106 81944 21582 82090
rect 21750 81944 22318 82090
rect 22486 81944 22962 82090
rect 23130 81944 23698 82090
rect 23866 81944 24342 82090
rect 24510 81944 25078 82090
rect 25246 81944 25722 82090
rect 25890 81944 26458 82090
rect 26626 81944 27102 82090
rect 27270 81944 27838 82090
rect 28006 81944 28482 82090
rect 28650 81944 29218 82090
rect 29386 81944 29862 82090
rect 30030 81944 30598 82090
rect 30766 81944 31242 82090
rect 31410 81944 31978 82090
rect 32146 81944 32622 82090
rect 32790 81944 33358 82090
rect 33526 81944 34002 82090
rect 34170 81944 34738 82090
rect 34906 81944 35382 82090
rect 35550 81944 36118 82090
rect 36286 81944 36762 82090
rect 36930 81944 37498 82090
rect 37666 81944 38234 82090
rect 38402 81944 38878 82090
rect 39046 81944 39614 82090
rect 39782 81944 40258 82090
rect 40426 81944 40994 82090
rect 41162 81944 41638 82090
rect 41806 81944 42374 82090
rect 42542 81944 43018 82090
rect 43186 81944 43754 82090
rect 43922 81944 44398 82090
rect 44566 81944 45134 82090
rect 45302 81944 45778 82090
rect 45946 81944 46514 82090
rect 46682 81944 47158 82090
rect 47326 81944 47894 82090
rect 48062 81944 48538 82090
rect 48706 81944 49274 82090
rect 49442 81944 49918 82090
rect 50086 81944 50654 82090
rect 50822 81944 51298 82090
rect 51466 81944 52034 82090
rect 52202 81944 52678 82090
rect 52846 81944 53414 82090
rect 53582 81944 54058 82090
rect 54226 81944 54794 82090
rect 54962 81944 55438 82090
rect 55606 81944 56174 82090
rect 56342 81944 56818 82090
rect 56986 81944 57554 82090
rect 57722 81944 58198 82090
rect 58366 81944 58934 82090
rect 59102 81944 59578 82090
rect 59746 81944 60314 82090
rect 60482 81944 60958 82090
rect 61126 81944 61694 82090
rect 61862 81944 62338 82090
rect 62506 81944 63074 82090
rect 63242 81944 63718 82090
rect 63886 81944 64454 82090
rect 64622 81944 65098 82090
rect 65266 81944 65834 82090
rect 66002 81944 66478 82090
rect 66646 81944 67214 82090
rect 67382 81944 67858 82090
rect 68026 81944 68594 82090
rect 68762 81944 69238 82090
rect 69406 81944 69974 82090
rect 70142 81944 70618 82090
rect 70786 81944 71354 82090
rect 71522 81944 71998 82090
rect 72166 81944 72734 82090
rect 72902 81944 73378 82090
rect 73546 81944 74114 82090
rect 74282 81944 74758 82090
rect 74926 81944 75494 82090
rect 75662 81944 75974 82090
rect 20 856 75974 81944
rect 20 2 146 856
rect 314 2 514 856
rect 682 2 882 856
rect 1050 2 1342 856
rect 1510 2 1710 856
rect 1878 2 2170 856
rect 2338 2 2538 856
rect 2706 2 2998 856
rect 3166 2 3366 856
rect 3534 2 3734 856
rect 3902 2 4194 856
rect 4362 2 4562 856
rect 4730 2 5022 856
rect 5190 2 5390 856
rect 5558 2 5850 856
rect 6018 2 6218 856
rect 6386 2 6678 856
rect 6846 2 7046 856
rect 7214 2 7414 856
rect 7582 2 7874 856
rect 8042 2 8242 856
rect 8410 2 8702 856
rect 8870 2 9070 856
rect 9238 2 9530 856
rect 9698 2 9898 856
rect 10066 2 10358 856
rect 10526 2 10726 856
rect 10894 2 11094 856
rect 11262 2 11554 856
rect 11722 2 11922 856
rect 12090 2 12382 856
rect 12550 2 12750 856
rect 12918 2 13210 856
rect 13378 2 13578 856
rect 13746 2 13946 856
rect 14114 2 14406 856
rect 14574 2 14774 856
rect 14942 2 15234 856
rect 15402 2 15602 856
rect 15770 2 16062 856
rect 16230 2 16430 856
rect 16598 2 16890 856
rect 17058 2 17258 856
rect 17426 2 17626 856
rect 17794 2 18086 856
rect 18254 2 18454 856
rect 18622 2 18914 856
rect 19082 2 19282 856
rect 19450 2 19742 856
rect 19910 2 20110 856
rect 20278 2 20570 856
rect 20738 2 20938 856
rect 21106 2 21306 856
rect 21474 2 21766 856
rect 21934 2 22134 856
rect 22302 2 22594 856
rect 22762 2 22962 856
rect 23130 2 23422 856
rect 23590 2 23790 856
rect 23958 2 24250 856
rect 24418 2 24618 856
rect 24786 2 24986 856
rect 25154 2 25446 856
rect 25614 2 25814 856
rect 25982 2 26274 856
rect 26442 2 26642 856
rect 26810 2 27102 856
rect 27270 2 27470 856
rect 27638 2 27838 856
rect 28006 2 28298 856
rect 28466 2 28666 856
rect 28834 2 29126 856
rect 29294 2 29494 856
rect 29662 2 29954 856
rect 30122 2 30322 856
rect 30490 2 30782 856
rect 30950 2 31150 856
rect 31318 2 31518 856
rect 31686 2 31978 856
rect 32146 2 32346 856
rect 32514 2 32806 856
rect 32974 2 33174 856
rect 33342 2 33634 856
rect 33802 2 34002 856
rect 34170 2 34462 856
rect 34630 2 34830 856
rect 34998 2 35198 856
rect 35366 2 35658 856
rect 35826 2 36026 856
rect 36194 2 36486 856
rect 36654 2 36854 856
rect 37022 2 37314 856
rect 37482 2 37682 856
rect 37850 2 38142 856
rect 38310 2 38510 856
rect 38678 2 38878 856
rect 39046 2 39338 856
rect 39506 2 39706 856
rect 39874 2 40166 856
rect 40334 2 40534 856
rect 40702 2 40994 856
rect 41162 2 41362 856
rect 41530 2 41730 856
rect 41898 2 42190 856
rect 42358 2 42558 856
rect 42726 2 43018 856
rect 43186 2 43386 856
rect 43554 2 43846 856
rect 44014 2 44214 856
rect 44382 2 44674 856
rect 44842 2 45042 856
rect 45210 2 45410 856
rect 45578 2 45870 856
rect 46038 2 46238 856
rect 46406 2 46698 856
rect 46866 2 47066 856
rect 47234 2 47526 856
rect 47694 2 47894 856
rect 48062 2 48354 856
rect 48522 2 48722 856
rect 48890 2 49090 856
rect 49258 2 49550 856
rect 49718 2 49918 856
rect 50086 2 50378 856
rect 50546 2 50746 856
rect 50914 2 51206 856
rect 51374 2 51574 856
rect 51742 2 51942 856
rect 52110 2 52402 856
rect 52570 2 52770 856
rect 52938 2 53230 856
rect 53398 2 53598 856
rect 53766 2 54058 856
rect 54226 2 54426 856
rect 54594 2 54886 856
rect 55054 2 55254 856
rect 55422 2 55622 856
rect 55790 2 56082 856
rect 56250 2 56450 856
rect 56618 2 56910 856
rect 57078 2 57278 856
rect 57446 2 57738 856
rect 57906 2 58106 856
rect 58274 2 58566 856
rect 58734 2 58934 856
rect 59102 2 59302 856
rect 59470 2 59762 856
rect 59930 2 60130 856
rect 60298 2 60590 856
rect 60758 2 60958 856
rect 61126 2 61418 856
rect 61586 2 61786 856
rect 61954 2 62246 856
rect 62414 2 62614 856
rect 62782 2 62982 856
rect 63150 2 63442 856
rect 63610 2 63810 856
rect 63978 2 64270 856
rect 64438 2 64638 856
rect 64806 2 65098 856
rect 65266 2 65466 856
rect 65634 2 65834 856
rect 66002 2 66294 856
rect 66462 2 66662 856
rect 66830 2 67122 856
rect 67290 2 67490 856
rect 67658 2 67950 856
rect 68118 2 68318 856
rect 68486 2 68778 856
rect 68946 2 69146 856
rect 69314 2 69514 856
rect 69682 2 69974 856
rect 70142 2 70342 856
rect 70510 2 70802 856
rect 70970 2 71170 856
rect 71338 2 71630 856
rect 71798 2 71998 856
rect 72166 2 72458 856
rect 72626 2 72826 856
rect 72994 2 73194 856
rect 73362 2 73654 856
rect 73822 2 74022 856
rect 74190 2 74482 856
rect 74650 2 74850 856
rect 75018 2 75310 856
rect 75478 2 75678 856
rect 75846 2 75974 856
<< metal3 >>
rect 75200 81744 76000 81864
rect 75200 79840 76000 79960
rect 0 78072 800 78192
rect 75200 77936 76000 78056
rect 75200 76032 76000 76152
rect 75200 74128 76000 74248
rect 75200 72224 76000 72344
rect 75200 70456 76000 70576
rect 0 68824 800 68944
rect 75200 68552 76000 68672
rect 75200 66648 76000 66768
rect 75200 64744 76000 64864
rect 75200 62840 76000 62960
rect 75200 60936 76000 61056
rect 0 59712 800 59832
rect 75200 59168 76000 59288
rect 75200 57264 76000 57384
rect 75200 55360 76000 55480
rect 75200 53456 76000 53576
rect 75200 51552 76000 51672
rect 0 50464 800 50584
rect 75200 49648 76000 49768
rect 75200 47880 76000 48000
rect 75200 45976 76000 46096
rect 75200 44072 76000 44192
rect 75200 42168 76000 42288
rect 0 41216 800 41336
rect 75200 40264 76000 40384
rect 75200 38360 76000 38480
rect 75200 36456 76000 36576
rect 75200 34688 76000 34808
rect 75200 32784 76000 32904
rect 0 32104 800 32224
rect 75200 30880 76000 31000
rect 75200 28976 76000 29096
rect 75200 27072 76000 27192
rect 75200 25168 76000 25288
rect 75200 23400 76000 23520
rect 0 22856 800 22976
rect 75200 21496 76000 21616
rect 75200 19592 76000 19712
rect 75200 17688 76000 17808
rect 75200 15784 76000 15904
rect 75200 13880 76000 14000
rect 0 13608 800 13728
rect 75200 12112 76000 12232
rect 75200 10208 76000 10328
rect 75200 8304 76000 8424
rect 75200 6400 76000 6520
rect 0 4496 800 4616
rect 75200 4496 76000 4616
rect 75200 2592 76000 2712
rect 75200 824 76000 944
<< obsm3 >>
rect 800 81664 75120 81837
rect 800 80040 75979 81664
rect 800 79760 75120 80040
rect 800 78272 75979 79760
rect 880 78136 75979 78272
rect 880 77992 75120 78136
rect 800 77856 75120 77992
rect 800 76232 75979 77856
rect 800 75952 75120 76232
rect 800 74328 75979 75952
rect 800 74048 75120 74328
rect 800 72424 75979 74048
rect 800 72144 75120 72424
rect 800 70656 75979 72144
rect 800 70376 75120 70656
rect 800 69024 75979 70376
rect 880 68752 75979 69024
rect 880 68744 75120 68752
rect 800 68472 75120 68744
rect 800 66848 75979 68472
rect 800 66568 75120 66848
rect 800 64944 75979 66568
rect 800 64664 75120 64944
rect 800 63040 75979 64664
rect 800 62760 75120 63040
rect 800 61136 75979 62760
rect 800 60856 75120 61136
rect 800 59912 75979 60856
rect 880 59632 75979 59912
rect 800 59368 75979 59632
rect 800 59088 75120 59368
rect 800 57464 75979 59088
rect 800 57184 75120 57464
rect 800 55560 75979 57184
rect 800 55280 75120 55560
rect 800 53656 75979 55280
rect 800 53376 75120 53656
rect 800 51752 75979 53376
rect 800 51472 75120 51752
rect 800 50664 75979 51472
rect 880 50384 75979 50664
rect 800 49848 75979 50384
rect 800 49568 75120 49848
rect 800 48080 75979 49568
rect 800 47800 75120 48080
rect 800 46176 75979 47800
rect 800 45896 75120 46176
rect 800 44272 75979 45896
rect 800 43992 75120 44272
rect 800 42368 75979 43992
rect 800 42088 75120 42368
rect 800 41416 75979 42088
rect 880 41136 75979 41416
rect 800 40464 75979 41136
rect 800 40184 75120 40464
rect 800 38560 75979 40184
rect 800 38280 75120 38560
rect 800 36656 75979 38280
rect 800 36376 75120 36656
rect 800 34888 75979 36376
rect 800 34608 75120 34888
rect 800 32984 75979 34608
rect 800 32704 75120 32984
rect 800 32304 75979 32704
rect 880 32024 75979 32304
rect 800 31080 75979 32024
rect 800 30800 75120 31080
rect 800 29176 75979 30800
rect 800 28896 75120 29176
rect 800 27272 75979 28896
rect 800 26992 75120 27272
rect 800 25368 75979 26992
rect 800 25088 75120 25368
rect 800 23600 75979 25088
rect 800 23320 75120 23600
rect 800 23056 75979 23320
rect 880 22776 75979 23056
rect 800 21696 75979 22776
rect 800 21416 75120 21696
rect 800 19792 75979 21416
rect 800 19512 75120 19792
rect 800 17888 75979 19512
rect 800 17608 75120 17888
rect 800 15984 75979 17608
rect 800 15704 75120 15984
rect 800 14080 75979 15704
rect 800 13808 75120 14080
rect 880 13800 75120 13808
rect 880 13528 75979 13800
rect 800 12312 75979 13528
rect 800 12032 75120 12312
rect 800 10408 75979 12032
rect 800 10128 75120 10408
rect 800 8504 75979 10128
rect 800 8224 75120 8504
rect 800 6600 75979 8224
rect 800 6320 75120 6600
rect 800 4696 75979 6320
rect 880 4416 75120 4696
rect 800 2792 75979 4416
rect 800 2512 75120 2792
rect 800 1024 75979 2512
rect 800 744 75120 1024
rect 800 35 75979 744
<< metal4 >>
rect 4208 2128 4528 80560
rect 19568 2128 19888 80560
rect 34928 2128 35248 80560
rect 50288 2128 50608 80560
rect 65648 2128 65968 80560
<< obsm4 >>
rect 1715 80640 75933 80749
rect 1715 2048 4128 80640
rect 4608 2048 19488 80640
rect 19968 2048 34848 80640
rect 35328 2048 50208 80640
rect 50688 2048 65568 80640
rect 66048 2048 75933 80640
rect 1715 35 75933 2048
<< labels >>
rlabel metal2 s 23018 82000 23074 82800 6 addrA0[0]
port 1 nsew signal output
rlabel metal3 s 0 59712 800 59832 6 addrA0[1]
port 2 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 addrA0[2]
port 3 nsew signal output
rlabel metal3 s 0 41216 800 41336 6 addrA0[3]
port 4 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 addrA0[4]
port 5 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 addrA0[5]
port 6 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 addrA0[6]
port 7 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 addrA0[7]
port 8 nsew signal output
rlabel metal2 s 22374 82000 22430 82800 6 addrA1[0]
port 9 nsew signal output
rlabel metal2 s 74814 82000 74870 82800 6 addrA1[1]
port 10 nsew signal output
rlabel metal2 s 74170 82000 74226 82800 6 addrA1[2]
port 11 nsew signal output
rlabel metal2 s 73434 82000 73490 82800 6 addrA1[3]
port 12 nsew signal output
rlabel metal2 s 72790 82000 72846 82800 6 addrA1[4]
port 13 nsew signal output
rlabel metal2 s 70674 82000 70730 82800 6 addrA1[5]
port 14 nsew signal output
rlabel metal2 s 71410 82000 71466 82800 6 addrA1[6]
port 15 nsew signal output
rlabel metal2 s 72054 82000 72110 82800 6 addrA1[7]
port 16 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 addrB0[0]
port 17 nsew signal output
rlabel metal3 s 75200 77936 76000 78056 6 addrB0[1]
port 18 nsew signal output
rlabel metal3 s 75200 76032 76000 76152 6 addrB0[2]
port 19 nsew signal output
rlabel metal3 s 75200 74128 76000 74248 6 addrB0[3]
port 20 nsew signal output
rlabel metal3 s 75200 72224 76000 72344 6 addrB0[4]
port 21 nsew signal output
rlabel metal3 s 75200 70456 76000 70576 6 addrB0[5]
port 22 nsew signal output
rlabel metal3 s 75200 68552 76000 68672 6 addrB0[6]
port 23 nsew signal output
rlabel metal3 s 75200 66648 76000 66768 6 addrB0[7]
port 24 nsew signal output
rlabel metal3 s 75200 64744 76000 64864 6 addrB0[8]
port 25 nsew signal output
rlabel metal3 s 75200 2592 76000 2712 6 addrB1[0]
port 26 nsew signal output
rlabel metal3 s 75200 824 76000 944 6 addrB1[1]
port 27 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 addrB1[2]
port 28 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 addrB1[3]
port 29 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 addrB1[4]
port 30 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 addrB1[5]
port 31 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 addrB1[6]
port 32 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 addrB1[7]
port 33 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 addrB1[8]
port 34 nsew signal output
rlabel metal3 s 0 78072 800 78192 6 csbA0
port 35 nsew signal output
rlabel metal2 s 75550 82000 75606 82800 6 csbA1
port 36 nsew signal output
rlabel metal3 s 75200 81744 76000 81864 6 csbB0
port 37 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 csbB1
port 38 nsew signal output
rlabel metal2 s 26514 82000 26570 82800 6 dinA0[0]
port 39 nsew signal output
rlabel metal2 s 33414 82000 33470 82800 6 dinA0[10]
port 40 nsew signal output
rlabel metal2 s 34058 82000 34114 82800 6 dinA0[11]
port 41 nsew signal output
rlabel metal2 s 34794 82000 34850 82800 6 dinA0[12]
port 42 nsew signal output
rlabel metal2 s 35438 82000 35494 82800 6 dinA0[13]
port 43 nsew signal output
rlabel metal2 s 36174 82000 36230 82800 6 dinA0[14]
port 44 nsew signal output
rlabel metal2 s 36818 82000 36874 82800 6 dinA0[15]
port 45 nsew signal output
rlabel metal2 s 37554 82000 37610 82800 6 dinA0[16]
port 46 nsew signal output
rlabel metal2 s 38290 82000 38346 82800 6 dinA0[17]
port 47 nsew signal output
rlabel metal2 s 38934 82000 38990 82800 6 dinA0[18]
port 48 nsew signal output
rlabel metal2 s 39670 82000 39726 82800 6 dinA0[19]
port 49 nsew signal output
rlabel metal2 s 27158 82000 27214 82800 6 dinA0[1]
port 50 nsew signal output
rlabel metal2 s 40314 82000 40370 82800 6 dinA0[20]
port 51 nsew signal output
rlabel metal2 s 41050 82000 41106 82800 6 dinA0[21]
port 52 nsew signal output
rlabel metal2 s 41694 82000 41750 82800 6 dinA0[22]
port 53 nsew signal output
rlabel metal2 s 42430 82000 42486 82800 6 dinA0[23]
port 54 nsew signal output
rlabel metal2 s 43074 82000 43130 82800 6 dinA0[24]
port 55 nsew signal output
rlabel metal2 s 43810 82000 43866 82800 6 dinA0[25]
port 56 nsew signal output
rlabel metal2 s 44454 82000 44510 82800 6 dinA0[26]
port 57 nsew signal output
rlabel metal2 s 45190 82000 45246 82800 6 dinA0[27]
port 58 nsew signal output
rlabel metal2 s 45834 82000 45890 82800 6 dinA0[28]
port 59 nsew signal output
rlabel metal2 s 46570 82000 46626 82800 6 dinA0[29]
port 60 nsew signal output
rlabel metal2 s 27894 82000 27950 82800 6 dinA0[2]
port 61 nsew signal output
rlabel metal2 s 47214 82000 47270 82800 6 dinA0[30]
port 62 nsew signal output
rlabel metal2 s 47950 82000 48006 82800 6 dinA0[31]
port 63 nsew signal output
rlabel metal2 s 28538 82000 28594 82800 6 dinA0[3]
port 64 nsew signal output
rlabel metal2 s 29274 82000 29330 82800 6 dinA0[4]
port 65 nsew signal output
rlabel metal2 s 29918 82000 29974 82800 6 dinA0[5]
port 66 nsew signal output
rlabel metal2 s 30654 82000 30710 82800 6 dinA0[6]
port 67 nsew signal output
rlabel metal2 s 31298 82000 31354 82800 6 dinA0[7]
port 68 nsew signal output
rlabel metal2 s 32034 82000 32090 82800 6 dinA0[8]
port 69 nsew signal output
rlabel metal2 s 32678 82000 32734 82800 6 dinA0[9]
port 70 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 dinB0[0]
port 71 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 dinB0[10]
port 72 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 dinB0[11]
port 73 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 dinB0[12]
port 74 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 dinB0[13]
port 75 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 dinB0[14]
port 76 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 dinB0[15]
port 77 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 dinB0[16]
port 78 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 dinB0[17]
port 79 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 dinB0[18]
port 80 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 dinB0[19]
port 81 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 dinB0[1]
port 82 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 dinB0[20]
port 83 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 dinB0[21]
port 84 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 dinB0[22]
port 85 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 dinB0[23]
port 86 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 dinB0[24]
port 87 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 dinB0[25]
port 88 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 dinB0[26]
port 89 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 dinB0[27]
port 90 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 dinB0[28]
port 91 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 dinB0[29]
port 92 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 dinB0[2]
port 93 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 dinB0[30]
port 94 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 dinB0[31]
port 95 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 dinB0[3]
port 96 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 dinB0[4]
port 97 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 dinB0[5]
port 98 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 dinB0[6]
port 99 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 dinB0[7]
port 100 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 dinB0[8]
port 101 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 dinB0[9]
port 102 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 sram12_dout0[0]
port 103 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 sram12_dout0[10]
port 104 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 sram12_dout0[11]
port 105 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 sram12_dout0[12]
port 106 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 sram12_dout0[13]
port 107 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 sram12_dout0[14]
port 108 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 sram12_dout0[15]
port 109 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 sram12_dout0[16]
port 110 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 sram12_dout0[17]
port 111 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 sram12_dout0[18]
port 112 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 sram12_dout0[19]
port 113 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 sram12_dout0[1]
port 114 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 sram12_dout0[20]
port 115 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 sram12_dout0[21]
port 116 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 sram12_dout0[22]
port 117 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 sram12_dout0[23]
port 118 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 sram12_dout0[24]
port 119 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 sram12_dout0[25]
port 120 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 sram12_dout0[26]
port 121 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 sram12_dout0[27]
port 122 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 sram12_dout0[28]
port 123 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 sram12_dout0[29]
port 124 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 sram12_dout0[2]
port 125 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 sram12_dout0[30]
port 126 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 sram12_dout0[31]
port 127 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 sram12_dout0[3]
port 128 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 sram12_dout0[4]
port 129 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 sram12_dout0[5]
port 130 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 sram12_dout0[6]
port 131 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 sram12_dout0[7]
port 132 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 sram12_dout0[8]
port 133 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 sram12_dout0[9]
port 134 nsew signal input
rlabel metal3 s 75200 4496 76000 4616 6 sram12_dout1[0]
port 135 nsew signal input
rlabel metal3 s 75200 23400 76000 23520 6 sram12_dout1[10]
port 136 nsew signal input
rlabel metal3 s 75200 25168 76000 25288 6 sram12_dout1[11]
port 137 nsew signal input
rlabel metal3 s 75200 27072 76000 27192 6 sram12_dout1[12]
port 138 nsew signal input
rlabel metal3 s 75200 28976 76000 29096 6 sram12_dout1[13]
port 139 nsew signal input
rlabel metal3 s 75200 30880 76000 31000 6 sram12_dout1[14]
port 140 nsew signal input
rlabel metal3 s 75200 32784 76000 32904 6 sram12_dout1[15]
port 141 nsew signal input
rlabel metal3 s 75200 34688 76000 34808 6 sram12_dout1[16]
port 142 nsew signal input
rlabel metal3 s 75200 36456 76000 36576 6 sram12_dout1[17]
port 143 nsew signal input
rlabel metal3 s 75200 38360 76000 38480 6 sram12_dout1[18]
port 144 nsew signal input
rlabel metal3 s 75200 40264 76000 40384 6 sram12_dout1[19]
port 145 nsew signal input
rlabel metal3 s 75200 6400 76000 6520 6 sram12_dout1[1]
port 146 nsew signal input
rlabel metal3 s 75200 42168 76000 42288 6 sram12_dout1[20]
port 147 nsew signal input
rlabel metal3 s 75200 44072 76000 44192 6 sram12_dout1[21]
port 148 nsew signal input
rlabel metal3 s 75200 45976 76000 46096 6 sram12_dout1[22]
port 149 nsew signal input
rlabel metal3 s 75200 47880 76000 48000 6 sram12_dout1[23]
port 150 nsew signal input
rlabel metal3 s 75200 49648 76000 49768 6 sram12_dout1[24]
port 151 nsew signal input
rlabel metal3 s 75200 51552 76000 51672 6 sram12_dout1[25]
port 152 nsew signal input
rlabel metal3 s 75200 53456 76000 53576 6 sram12_dout1[26]
port 153 nsew signal input
rlabel metal3 s 75200 55360 76000 55480 6 sram12_dout1[27]
port 154 nsew signal input
rlabel metal3 s 75200 57264 76000 57384 6 sram12_dout1[28]
port 155 nsew signal input
rlabel metal3 s 75200 59168 76000 59288 6 sram12_dout1[29]
port 156 nsew signal input
rlabel metal3 s 75200 8304 76000 8424 6 sram12_dout1[2]
port 157 nsew signal input
rlabel metal3 s 75200 60936 76000 61056 6 sram12_dout1[30]
port 158 nsew signal input
rlabel metal3 s 75200 62840 76000 62960 6 sram12_dout1[31]
port 159 nsew signal input
rlabel metal3 s 75200 10208 76000 10328 6 sram12_dout1[3]
port 160 nsew signal input
rlabel metal3 s 75200 12112 76000 12232 6 sram12_dout1[4]
port 161 nsew signal input
rlabel metal3 s 75200 13880 76000 14000 6 sram12_dout1[5]
port 162 nsew signal input
rlabel metal3 s 75200 15784 76000 15904 6 sram12_dout1[6]
port 163 nsew signal input
rlabel metal3 s 75200 17688 76000 17808 6 sram12_dout1[7]
port 164 nsew signal input
rlabel metal3 s 75200 19592 76000 19712 6 sram12_dout1[8]
port 165 nsew signal input
rlabel metal3 s 75200 21496 76000 21616 6 sram12_dout1[9]
port 166 nsew signal input
rlabel metal2 s 48594 82000 48650 82800 6 sram1_dout0[0]
port 167 nsew signal input
rlabel metal2 s 55494 82000 55550 82800 6 sram1_dout0[10]
port 168 nsew signal input
rlabel metal2 s 56230 82000 56286 82800 6 sram1_dout0[11]
port 169 nsew signal input
rlabel metal2 s 56874 82000 56930 82800 6 sram1_dout0[12]
port 170 nsew signal input
rlabel metal2 s 57610 82000 57666 82800 6 sram1_dout0[13]
port 171 nsew signal input
rlabel metal2 s 58254 82000 58310 82800 6 sram1_dout0[14]
port 172 nsew signal input
rlabel metal2 s 58990 82000 59046 82800 6 sram1_dout0[15]
port 173 nsew signal input
rlabel metal2 s 59634 82000 59690 82800 6 sram1_dout0[16]
port 174 nsew signal input
rlabel metal2 s 60370 82000 60426 82800 6 sram1_dout0[17]
port 175 nsew signal input
rlabel metal2 s 61014 82000 61070 82800 6 sram1_dout0[18]
port 176 nsew signal input
rlabel metal2 s 61750 82000 61806 82800 6 sram1_dout0[19]
port 177 nsew signal input
rlabel metal2 s 49330 82000 49386 82800 6 sram1_dout0[1]
port 178 nsew signal input
rlabel metal2 s 62394 82000 62450 82800 6 sram1_dout0[20]
port 179 nsew signal input
rlabel metal2 s 63130 82000 63186 82800 6 sram1_dout0[21]
port 180 nsew signal input
rlabel metal2 s 63774 82000 63830 82800 6 sram1_dout0[22]
port 181 nsew signal input
rlabel metal2 s 64510 82000 64566 82800 6 sram1_dout0[23]
port 182 nsew signal input
rlabel metal2 s 65154 82000 65210 82800 6 sram1_dout0[24]
port 183 nsew signal input
rlabel metal2 s 65890 82000 65946 82800 6 sram1_dout0[25]
port 184 nsew signal input
rlabel metal2 s 66534 82000 66590 82800 6 sram1_dout0[26]
port 185 nsew signal input
rlabel metal2 s 67270 82000 67326 82800 6 sram1_dout0[27]
port 186 nsew signal input
rlabel metal2 s 67914 82000 67970 82800 6 sram1_dout0[28]
port 187 nsew signal input
rlabel metal2 s 68650 82000 68706 82800 6 sram1_dout0[29]
port 188 nsew signal input
rlabel metal2 s 49974 82000 50030 82800 6 sram1_dout0[2]
port 189 nsew signal input
rlabel metal2 s 69294 82000 69350 82800 6 sram1_dout0[30]
port 190 nsew signal input
rlabel metal2 s 70030 82000 70086 82800 6 sram1_dout0[31]
port 191 nsew signal input
rlabel metal2 s 50710 82000 50766 82800 6 sram1_dout0[3]
port 192 nsew signal input
rlabel metal2 s 51354 82000 51410 82800 6 sram1_dout0[4]
port 193 nsew signal input
rlabel metal2 s 52090 82000 52146 82800 6 sram1_dout0[5]
port 194 nsew signal input
rlabel metal2 s 52734 82000 52790 82800 6 sram1_dout0[6]
port 195 nsew signal input
rlabel metal2 s 53470 82000 53526 82800 6 sram1_dout0[7]
port 196 nsew signal input
rlabel metal2 s 54114 82000 54170 82800 6 sram1_dout0[8]
port 197 nsew signal input
rlabel metal2 s 54850 82000 54906 82800 6 sram1_dout0[9]
port 198 nsew signal input
rlabel metal2 s 294 82000 350 82800 6 sram1_dout1[0]
port 199 nsew signal input
rlabel metal2 s 7194 82000 7250 82800 6 sram1_dout1[10]
port 200 nsew signal input
rlabel metal2 s 7838 82000 7894 82800 6 sram1_dout1[11]
port 201 nsew signal input
rlabel metal2 s 8574 82000 8630 82800 6 sram1_dout1[12]
port 202 nsew signal input
rlabel metal2 s 9218 82000 9274 82800 6 sram1_dout1[13]
port 203 nsew signal input
rlabel metal2 s 9954 82000 10010 82800 6 sram1_dout1[14]
port 204 nsew signal input
rlabel metal2 s 10598 82000 10654 82800 6 sram1_dout1[15]
port 205 nsew signal input
rlabel metal2 s 11334 82000 11390 82800 6 sram1_dout1[16]
port 206 nsew signal input
rlabel metal2 s 11978 82000 12034 82800 6 sram1_dout1[17]
port 207 nsew signal input
rlabel metal2 s 12714 82000 12770 82800 6 sram1_dout1[18]
port 208 nsew signal input
rlabel metal2 s 13358 82000 13414 82800 6 sram1_dout1[19]
port 209 nsew signal input
rlabel metal2 s 938 82000 994 82800 6 sram1_dout1[1]
port 210 nsew signal input
rlabel metal2 s 14094 82000 14150 82800 6 sram1_dout1[20]
port 211 nsew signal input
rlabel metal2 s 14738 82000 14794 82800 6 sram1_dout1[21]
port 212 nsew signal input
rlabel metal2 s 15474 82000 15530 82800 6 sram1_dout1[22]
port 213 nsew signal input
rlabel metal2 s 16118 82000 16174 82800 6 sram1_dout1[23]
port 214 nsew signal input
rlabel metal2 s 16854 82000 16910 82800 6 sram1_dout1[24]
port 215 nsew signal input
rlabel metal2 s 17498 82000 17554 82800 6 sram1_dout1[25]
port 216 nsew signal input
rlabel metal2 s 18234 82000 18290 82800 6 sram1_dout1[26]
port 217 nsew signal input
rlabel metal2 s 18878 82000 18934 82800 6 sram1_dout1[27]
port 218 nsew signal input
rlabel metal2 s 19614 82000 19670 82800 6 sram1_dout1[28]
port 219 nsew signal input
rlabel metal2 s 20258 82000 20314 82800 6 sram1_dout1[29]
port 220 nsew signal input
rlabel metal2 s 1674 82000 1730 82800 6 sram1_dout1[2]
port 221 nsew signal input
rlabel metal2 s 20994 82000 21050 82800 6 sram1_dout1[30]
port 222 nsew signal input
rlabel metal2 s 21638 82000 21694 82800 6 sram1_dout1[31]
port 223 nsew signal input
rlabel metal2 s 2318 82000 2374 82800 6 sram1_dout1[3]
port 224 nsew signal input
rlabel metal2 s 3054 82000 3110 82800 6 sram1_dout1[4]
port 225 nsew signal input
rlabel metal2 s 3698 82000 3754 82800 6 sram1_dout1[5]
port 226 nsew signal input
rlabel metal2 s 4434 82000 4490 82800 6 sram1_dout1[6]
port 227 nsew signal input
rlabel metal2 s 5078 82000 5134 82800 6 sram1_dout1[7]
port 228 nsew signal input
rlabel metal2 s 5814 82000 5870 82800 6 sram1_dout1[8]
port 229 nsew signal input
rlabel metal2 s 6458 82000 6514 82800 6 sram1_dout1[9]
port 230 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 user_irq[0]
port 231 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 user_irq[1]
port 232 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 user_irq[2]
port 233 nsew signal output
rlabel metal4 s 4208 2128 4528 80560 6 vccd1
port 234 nsew power input
rlabel metal4 s 34928 2128 35248 80560 6 vccd1
port 234 nsew power input
rlabel metal4 s 65648 2128 65968 80560 6 vccd1
port 234 nsew power input
rlabel metal4 s 19568 2128 19888 80560 6 vssd1
port 235 nsew ground input
rlabel metal4 s 50288 2128 50608 80560 6 vssd1
port 235 nsew ground input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 236 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 237 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_ack_o
port 238 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_adr_i[0]
port 239 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[10]
port 240 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[11]
port 241 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[12]
port 242 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[13]
port 243 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[14]
port 244 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_adr_i[15]
port 245 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[16]
port 246 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[17]
port 247 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[18]
port 248 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[19]
port 249 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[1]
port 250 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[20]
port 251 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[21]
port 252 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[22]
port 253 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[23]
port 254 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_adr_i[24]
port 255 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_adr_i[25]
port 256 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[26]
port 257 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[27]
port 258 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_adr_i[28]
port 259 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_adr_i[29]
port 260 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_adr_i[2]
port 261 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_adr_i[30]
port 262 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 wbs_adr_i[31]
port 263 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[3]
port 264 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[4]
port 265 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[5]
port 266 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_adr_i[6]
port 267 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_adr_i[7]
port 268 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[8]
port 269 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_adr_i[9]
port 270 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_cyc_i
port 271 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_dat_i[0]
port 272 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_i[10]
port 273 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[11]
port 274 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[12]
port 275 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[13]
port 276 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_i[14]
port 277 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[15]
port 278 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_i[16]
port 279 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_i[17]
port 280 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[18]
port 281 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_i[19]
port 282 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[1]
port 283 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_i[20]
port 284 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_i[21]
port 285 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wbs_dat_i[22]
port 286 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_i[23]
port 287 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_i[24]
port 288 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_i[25]
port 289 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_dat_i[26]
port 290 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_i[27]
port 291 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_i[28]
port 292 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[29]
port 293 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[2]
port 294 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_i[30]
port 295 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_dat_i[31]
port 296 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_i[3]
port 297 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[4]
port 298 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[5]
port 299 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_i[6]
port 300 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[7]
port 301 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_i[8]
port 302 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[9]
port 303 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_o[0]
port 304 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_o[10]
port 305 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[11]
port 306 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[12]
port 307 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[13]
port 308 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[14]
port 309 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_o[15]
port 310 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[16]
port 311 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_o[17]
port 312 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[18]
port 313 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_o[19]
port 314 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[1]
port 315 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[20]
port 316 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_o[21]
port 317 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[22]
port 318 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_o[23]
port 319 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_o[24]
port 320 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[25]
port 321 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[26]
port 322 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_o[27]
port 323 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_o[28]
port 324 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 wbs_dat_o[29]
port 325 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_o[2]
port 326 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_o[30]
port 327 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 wbs_dat_o[31]
port 328 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[3]
port 329 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[4]
port 330 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[5]
port 331 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[6]
port 332 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_o[7]
port 333 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[8]
port 334 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[9]
port 335 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[0]
port 336 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_sel_i[1]
port 337 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_sel_i[2]
port 338 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_sel_i[3]
port 339 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_stb_i
port 340 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_we_i
port 341 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 webA
port 342 nsew signal output
rlabel metal3 s 75200 79840 76000 79960 6 webB
port 343 nsew signal output
rlabel metal2 s 23754 82000 23810 82800 6 wmaskA[0]
port 344 nsew signal output
rlabel metal2 s 24398 82000 24454 82800 6 wmaskA[1]
port 345 nsew signal output
rlabel metal2 s 25134 82000 25190 82800 6 wmaskA[2]
port 346 nsew signal output
rlabel metal2 s 25778 82000 25834 82800 6 wmaskA[3]
port 347 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 wmaskB[0]
port 348 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 wmaskB[1]
port 349 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 wmaskB[2]
port 350 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 wmaskB[3]
port 351 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 76000 82800
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 21642862
string GDS_FILE /home/re19/Caravel/temporal_runtime_monitor/openlane/user_project/runs/user_project/results/finishing/user_project.magic.gds
string GDS_START 1461590
<< end >>

